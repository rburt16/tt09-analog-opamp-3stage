** sch_path: /foss/designs/tt09-analog-opamp-3stage/xschem/tb_op_amp_3stage.sch
**.subckt tb_op_amp_3stage
Vin in+ GND 0.9 AC 1 pulse 0.1 1.2 0 10n 10n 500n 1u
Vsupply VDPWR GND 1.8
Rload out net1 10k m=1
Vsupply1 net1 GND 0.9
Rload1 net2 net1 100 m=1
Cload out net1 1f m=1
Cload1 out net2 1f m=1
I7 x1.cmfb GND 0 pulse 0u 0u 0 2n 2n 500n 1u
x1 VDPWR out in- in+ GND op_amp_3stage
Rfeedback out in- 1 m=1
Vin1 net3 GND 0.9 pulse 0.1 1.7 0 10n 10n 500n 1u
Rfb2 GND net3 5k m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.control
.option savecurrents
*.options temp=125
dc Vin 0.1 1.2 0.02
*temp -40 125 15
plot v(in+) v(x1.commonmode) v(VDPWR)
plot v(out) v(x1.pdrive) v(x1.ndrive)
plot v(in+)-v(in-) ylimit 100u -100u ydelta 50u
plot @m.x1.xm2.msky130_fd_pr__pfet_01v8_lvt[id] @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
plot 1/(@m.x1.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]+@m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gm])
*plot i(Vmeas) title vs_Supply_tt_-40degto125deg
ac dec 100 1 1e9
plot db(v(out)/v(in+,in-)) ph(v(out)/v(in+,in-))*57.3 ylimit 180 -180 ydelta 20
plot db(v(out)/v(x1.in+2,x1.in-2)) ph(v(out)/v(x1.in+2,x1.in-2))*57.3 ylimit 180 -180 ydelta 20
plot db(v(out)) xlog ylimit 6 -6 ydelta 3
dc temp -40 125 5
*plot v(out) v(pdrive) v(ndrive)
*plot i(Vmeas) title vs_Temp_tt
*plot v(x1.drive) title vs_Temp_tt
*plot v(x1.ptat) title vs_Temp_tt
*set temp=-40
*tran 2n 1u
*plot v(VSS) title Start_Up_tt_-40deg
*plot v(x1.ptat) title Stability
*plot i(Vmeas) @m.x1.xm18.msky130_fd_pr__nfet_01v8[id] title Start_Up_tt
*set temp=125
tran 2n 1u
plot v(out) v(x1.pdrive) v(x1.ndrive)
plot @m.x1.xm2.msky130_fd_pr__pfet_01v8_lvt[id]
*plot v(out) ylimit 0.86 1.04 ydelta 0.02
plot v(out)
plot v(x1.cmfb)
*plot V(VSS) title Start_Up_tt_125deg
*plot v(x1.ptat)
*plot i(Vmeas) @m.x1.xm18.msky130_fd_pr__nfet_01v8[id] title Start_Up_tt_125deg
noise v(out) Vin dec 10 1 100MEG 1
write noise1.all noise2.all
setplot noise1
setplot noise2
plot onoise_spectrum xlog ylog
*plot onoise.m.x1.xm15.msky130_fd_pr__pfet_01v8_lvt onoise.m.x1.xm14.msky130_fd_pr__nfet_01v8_lvt xlog ylog
*plot onoise.m.x1.xm14.msky130_fd_pr__nfet_01v8_lvt onoise.m.x1.xm14.msky130_fd_pr__nfet_01v8_lvt.id xlog ylog
save all
*set temp=27
op
print all
write tb_op_amp_3stage.raw
.endc
.save all @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gm] @m.x1.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
+ @m.x1.xm11.msky130_fd_pr__pfet_01v8[gm] @m.x1.xm12.msky130_fd_pr__pfet_01v8[gm]
+ @m.x1.xm15.msky130_fd_pr__pfet_01v8_lvt[gm] @m.x1.xm16.msky130_fd_pr__pfet_01v8_lvt[gm]
+ @m.x1.xm14.msky130_fd_pr__nfet_01v8_lvt[gm] @m.x1.xm13.msky130_fd_pr__nfet_01v8_lvt[gm]


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/tt09-analog-opamp-3stage/xschem/op_amp_3stage.sym # of pins=5
** sym_path: /foss/designs/tt09-analog-opamp-3stage/xschem/op_amp_3stage.sym
** sch_path: /foss/designs/tt09-analog-opamp-3stage/xschem/op_amp_3stage.sch
.subckt op_amp_3stage VDPWR out in- in+ VGND
*.opin out
*.ipin VDPWR
*.ipin VGND
*.ipin in-
*.ipin in+
XM2 out pdrive VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=110 nf=11 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM6 net2 net2 VDPWR VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 ndrive I2_10uA<-- pdrive VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 I2_10uA<-- I2_10uA<-- net2 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 <--I3_10uA <--I3_10uA net1 VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 pdrive <--I3_10uA ndrive VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 out ndrive VGND VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=42.5 nf=17 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM9 ndrive net3 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=1.0 W=2.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net3 net3 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=1.0 W=2.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net3 in-2 <--I4_20uA VDPWR sky130_fd_pr__pfet_01v8 L=0.7 W=20 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 ndrive in+2 <--I4_20uA VDPWR sky130_fd_pr__pfet_01v8 L=0.7 W=20 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 out ndrive sky130_fd_pr__cap_mim_m3_1 W=27 L=10 MF=1 m=1
XC2 out pdrive sky130_fd_pr__cap_mim_m3_1 W=27 L=10 MF=1 m=1
XM13 in-2 net4 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=8 W=40 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 in+2 net4 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=8 W=40 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC3 VGND in+2 sky130_fd_pr__cap_mim_m3_1 W=109 L=30 MF=1 m=1
XC4 out in-2 sky130_fd_pr__cap_mim_m3_1 W=109 L=30 MF=1 m=1
XM15 in+2 in- commonmode VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.7 W=640 nf=32 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM16 in-2 in+ commonmode VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.7 W=640 nf=32 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM19 net4 net4 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=8 W=40 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 net4 VGND net5 VDPWR sky130_fd_pr__pfet_01v8 L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 VGND in+2 cmfb VDPWR sky130_fd_pr__pfet_01v8 L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 VGND in-2 cmfb VDPWR sky130_fd_pr__pfet_01v8 L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 VDPWR net6 VGND bias_generator
XM21 net6 net6 net7 VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM23 net9 net6 net8 VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=30 nf=10 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM25 net10 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM26 net11 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM27 net12 net9 net10 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM28 net9 net9 net11 VDPWR sky130_fd_pr__pfet_01v8_lvt L=.35 W=10.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM22 net7 net7 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM24 net8 net7 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
XM29 net12 net12 net13 VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM30 I2_10uA<-- net12 net14 VGND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM31 net13 net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM32 net14 net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM34 ndrive net13 VGND VGND sky130_fd_pr__nfet_01v8_lvt L=4.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM33 net15 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM35 <--I3_10uA net9 net15 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM36 net16 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM37 pdrive net9 net16 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM38 net17 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM39 <--I4_20uA net9 net17 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM40 net18 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM41 commonmode net9 net18 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM42 net19 net9 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=30 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM43 cmfb net9 net19 VDPWR sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM44 net5 VGND cmfb VDPWR sky130_fd_pr__pfet_01v8 L=0.35 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/tt09-analog-opamp-3stage/xschem/bias_generator.sym # of pins=3
** sym_path: /foss/designs/tt09-analog-opamp-3stage/xschem/bias_generator.sym
** sch_path: /foss/designs/tt09-analog-opamp-3stage/xschem/bias_generator.sch
.subckt bias_generator VDPWR i_out VGND
*.ipin VGND
*.ipin VDPWR
*.opin i_out
XM9 ncascode ncascode net1 VGND sky130_fd_pr__nfet_01v8_lvt L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 pgate ncascode net4 VGND sky130_fd_pr__nfet_01v8_lvt L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net4 net1 ptat VGND sky130_fd_pr__nfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XM18 pgate startup VGND VGND sky130_fd_pr__nfet_01v8 L=8.0 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 startup net1 VGND VGND sky130_fd_pr__nfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 ptat drive VGND VGND sky130_fd_pr__nfet_01v8 L=8.0 W=1.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM7 drive drive net3 VGND sky130_fd_pr__nfet_01v8 L=13.1 W=1.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net3 drive ptat VGND sky130_fd_pr__nfet_01v8 L=8.0 W=1.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 pgate VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net6 pgate VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net7 pgate VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net5 pgate VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 startup net1 VDPWR VDPWR sky130_fd_pr__pfet_01v8 L=8.0 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 pgate pgate net2 VDPWR sky130_fd_pr__pfet_01v8_lvt L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 drive pgate net6 VDPWR sky130_fd_pr__pfet_01v8_lvt L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 i_out pgate net7 VDPWR sky130_fd_pr__pfet_01v8_lvt L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 ncascode pgate net5 VDPWR sky130_fd_pr__pfet_01v8_lvt L=1.0 W=8.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
