magic
tech sky130A
magscale 1 2
timestamp 1730563144
<< nwell >>
rect -32020 27340 -32018 27420
rect -31590 27120 -31588 27198
rect -40780 17110 -40750 17270
<< metal1 >>
rect -30150 29550 -30070 29560
rect -41660 29510 -41480 29540
rect -40810 29520 -31900 29550
rect -30150 29520 -30140 29550
rect -41660 29160 -41630 29510
rect -31930 29490 -30140 29520
rect -30080 29490 -30070 29550
rect -40590 29480 -40510 29490
rect -40590 29440 -40580 29480
rect -41490 29420 -40580 29440
rect -40520 29440 -40510 29480
rect -40520 29420 -37520 29440
rect -41490 29410 -37520 29420
rect -37660 29280 -37580 29290
rect -37660 29240 -37650 29280
rect -41290 29210 -40150 29240
rect -41290 29050 -41260 29210
rect -40770 29050 -40740 29210
rect -40180 29050 -40150 29210
rect -40050 29220 -37650 29240
rect -37590 29220 -37580 29280
rect -40050 29210 -37580 29220
rect -40050 29050 -40010 29210
rect -37550 28120 -37520 29410
rect -32080 29390 -31080 29420
rect -30470 29390 -30360 29420
rect -37430 29280 -37350 29290
rect -37430 29220 -37420 29280
rect -37360 29220 -37350 29280
rect -37430 29210 -37350 29220
rect -32080 28410 -32050 29390
rect -31190 29000 -31160 29390
rect -30470 29030 -30440 29390
rect -31050 29000 -30430 29030
rect -30320 29000 -30290 29490
rect -30150 29480 -30070 29490
rect -32330 28400 -32250 28410
rect -32330 28340 -32320 28400
rect -32260 28360 -32250 28400
rect -32150 28400 -32050 28410
rect -32150 28360 -32140 28400
rect -32260 28340 -32140 28360
rect -32080 28340 -32050 28400
rect -32330 28330 -32050 28340
rect -35690 28270 -32110 28300
rect -35690 28260 -35610 28270
rect -35690 28200 -35680 28260
rect -35620 28200 -35610 28260
rect -35690 28190 -35610 28200
rect -37550 28090 -33810 28120
rect -36600 27860 -36520 27870
rect -36600 27820 -36590 27860
rect -37110 27800 -36590 27820
rect -36530 27800 -36520 27860
rect -37110 27790 -36520 27800
rect -37110 27740 -37080 27790
rect -36600 27740 -36570 27790
rect -41550 27620 -41520 27670
rect -41030 27620 -41000 27670
rect -41660 27590 -41000 27620
rect -41660 27210 -41630 27560
rect -40590 27350 -40510 27360
rect -40590 27310 -40580 27350
rect -41490 27290 -40580 27310
rect -40520 27310 -40510 27350
rect -40520 27290 -40080 27310
rect -41490 27280 -40080 27290
rect -39940 27210 -39910 27560
rect -41660 27180 -37460 27210
rect -41660 25460 -41630 27180
rect -39870 26920 -37750 26950
rect -40590 26790 -40510 26800
rect -40590 26750 -40580 26790
rect -41490 26730 -40580 26750
rect -40520 26750 -40510 26790
rect -40520 26740 -39900 26750
rect -40520 26730 -39970 26740
rect -41490 26720 -39970 26730
rect -40780 26480 -40700 26490
rect -40780 26440 -40770 26480
rect -41290 26420 -40770 26440
rect -40710 26420 -40700 26480
rect -41290 26410 -40700 26420
rect -41290 26360 -41260 26410
rect -40770 26360 -40740 26410
rect -41550 24920 -41520 24980
rect -41030 24920 -41000 24980
rect -41650 24890 -41000 24920
rect -40590 24620 -40560 26720
rect -39980 26680 -39970 26720
rect -39910 26680 -39900 26740
rect -39980 26670 -39900 26680
rect -40220 26480 -40140 26490
rect -40530 26450 -40450 26460
rect -40530 26390 -40520 26450
rect -40460 26390 -40450 26450
rect -40220 26420 -40210 26480
rect -40150 26420 -40140 26480
rect -40220 26410 -40140 26420
rect -40530 26380 -40450 26390
rect -41490 24590 -40780 24620
rect -40590 24610 -40510 24620
rect -41490 24580 -40700 24590
rect -41490 24520 -40770 24580
rect -40710 24520 -40700 24580
rect -41490 24510 -40700 24520
rect -40590 24550 -40580 24610
rect -40520 24550 -40510 24610
rect -40590 24540 -40510 24550
rect -41490 24480 -40780 24510
rect -40780 24240 -40700 24250
rect -40780 24200 -40770 24240
rect -41290 24180 -40770 24200
rect -40710 24180 -40700 24240
rect -41290 24170 -40700 24180
rect -41290 24120 -41260 24170
rect -40770 24120 -40740 24170
rect -41550 22680 -41520 22740
rect -41030 22680 -41000 22740
rect -41660 22650 -41000 22680
rect -40590 22390 -40560 24540
rect -40480 24280 -40450 26380
rect -40180 26360 -40150 26410
rect -39870 26360 -39840 26920
rect -39690 26770 -37990 26780
rect -39690 26710 -39680 26770
rect -39620 26750 -37990 26770
rect -39620 26710 -39610 26750
rect -39690 26700 -39610 26710
rect -38690 26510 -38610 26520
rect -38690 26470 -38680 26510
rect -39200 26450 -38680 26470
rect -38620 26450 -38610 26510
rect -39200 26440 -38610 26450
rect -39200 26390 -39170 26440
rect -38680 26390 -38650 26440
rect -40040 26330 -39840 26360
rect -40140 24590 -40080 24620
rect -40220 24580 -40080 24590
rect -40220 24520 -40210 24580
rect -40150 24520 -40080 24580
rect -40220 24510 -40080 24520
rect -40140 24480 -40080 24510
rect -40480 24270 -40400 24280
rect -40480 24210 -40470 24270
rect -40410 24210 -40400 24270
rect -40480 24200 -40400 24210
rect -40220 24240 -40140 24250
rect -40590 22380 -40510 22390
rect -41490 22360 -40780 22380
rect -41490 22350 -40700 22360
rect -41490 22290 -40770 22350
rect -40710 22290 -40700 22350
rect -41490 22280 -40700 22290
rect -40590 22320 -40580 22380
rect -40520 22320 -40510 22380
rect -40590 22310 -40510 22320
rect -41490 22250 -40780 22280
rect -40780 22020 -40700 22030
rect -40780 21980 -40770 22020
rect -41290 21960 -40770 21980
rect -40710 21960 -40700 22020
rect -41290 21950 -40700 21960
rect -41290 21890 -41260 21950
rect -40770 21890 -40740 21950
rect -41550 20450 -41520 20510
rect -41030 20450 -41000 20510
rect -41660 20420 -41000 20450
rect -40590 20150 -40560 22310
rect -40480 22060 -40450 24200
rect -40220 24180 -40210 24240
rect -40150 24180 -40140 24240
rect -40220 24170 -40140 24180
rect -40180 24120 -40150 24170
rect -40030 24090 -40000 25010
rect -39460 24960 -39430 25010
rect -38940 24960 -38910 25010
rect -39570 24930 -38910 24960
rect -38500 24650 -38470 26750
rect -38320 26540 -38240 26550
rect -38320 26480 -38310 26540
rect -38250 26480 -38240 26540
rect -38320 26470 -38240 26480
rect -39400 24620 -38690 24650
rect -38500 24640 -38420 24650
rect -39400 24610 -38610 24620
rect -39400 24550 -38680 24610
rect -38620 24550 -38610 24610
rect -39400 24540 -38610 24550
rect -38500 24580 -38490 24640
rect -38430 24580 -38420 24640
rect -38500 24570 -38420 24580
rect -39400 24510 -38690 24540
rect -38690 24270 -38610 24280
rect -38690 24230 -38680 24270
rect -39200 24210 -38680 24230
rect -38620 24210 -38610 24270
rect -39200 24200 -38610 24210
rect -39200 24150 -39170 24200
rect -38690 24150 -38660 24200
rect -40140 22360 -40080 22380
rect -40220 22350 -40080 22360
rect -40220 22290 -40210 22350
rect -40150 22290 -40080 22350
rect -40220 22280 -40080 22290
rect -40140 22240 -40080 22280
rect -40480 22050 -40400 22060
rect -40480 21990 -40470 22050
rect -40410 21990 -40400 22050
rect -40480 21980 -40400 21990
rect -40220 22020 -40140 22030
rect -41490 20120 -40780 20150
rect -40590 20140 -40510 20150
rect -41490 20110 -40700 20120
rect -41490 20050 -40770 20110
rect -40710 20050 -40700 20110
rect -41490 20040 -40700 20050
rect -40590 20080 -40580 20140
rect -40520 20080 -40510 20140
rect -40590 20070 -40510 20080
rect -41490 20010 -40780 20040
rect -40780 19770 -40700 19780
rect -40780 19730 -40770 19770
rect -41290 19710 -40770 19730
rect -40710 19710 -40700 19770
rect -41290 19700 -40700 19710
rect -41290 19650 -41260 19700
rect -40770 19650 -40740 19700
rect -41660 18210 -41630 19170
rect -41550 18210 -41520 18270
rect -41030 18210 -41000 18270
rect -41660 18180 -41000 18210
rect -41660 17810 -41630 18180
rect -40590 17990 -40560 20070
rect -40480 19810 -40450 21980
rect -40220 21960 -40210 22020
rect -40150 21960 -40140 22020
rect -40220 21950 -40140 21960
rect -40180 21890 -40150 21950
rect -40030 21850 -40000 22770
rect -39460 22720 -39430 22770
rect -38940 22720 -38910 22770
rect -39570 22690 -38910 22720
rect -38500 22410 -38470 24570
rect -38270 24310 -38240 26470
rect -38130 26510 -38050 26520
rect -38130 26450 -38120 26510
rect -38060 26450 -38050 26510
rect -38130 26440 -38050 26450
rect -38080 26390 -38050 26440
rect -37890 25610 -37810 25620
rect -37890 25570 -37880 25610
rect -37960 25550 -37880 25570
rect -37820 25550 -37810 25610
rect -37960 25540 -37810 25550
rect -38050 24620 -37980 24650
rect -38130 24610 -37980 24620
rect -38130 24550 -38120 24610
rect -38060 24550 -37980 24610
rect -38130 24540 -37980 24550
rect -38050 24510 -37980 24540
rect -38320 24300 -38240 24310
rect -38320 24240 -38310 24300
rect -38250 24240 -38240 24300
rect -38320 24230 -38240 24240
rect -39400 22380 -38690 22410
rect -38500 22400 -38420 22410
rect -39400 22370 -38610 22380
rect -39400 22310 -38680 22370
rect -38620 22310 -38610 22370
rect -39400 22300 -38610 22310
rect -38500 22340 -38490 22400
rect -38430 22340 -38420 22400
rect -38500 22330 -38420 22340
rect -39400 22270 -38690 22300
rect -38690 22040 -38610 22050
rect -38690 22000 -38680 22040
rect -39200 21980 -38680 22000
rect -38620 21980 -38610 22040
rect -39200 21970 -38610 21980
rect -39200 21920 -39170 21970
rect -38690 21920 -38660 21970
rect -40140 20120 -40080 20150
rect -40220 20110 -40080 20120
rect -40220 20050 -40210 20110
rect -40150 20050 -40080 20110
rect -40220 20040 -40080 20050
rect -40140 20010 -40080 20040
rect -40480 19800 -40400 19810
rect -40480 19740 -40470 19800
rect -40410 19740 -40400 19800
rect -40480 19730 -40400 19740
rect -40220 19770 -40140 19780
rect -40220 19710 -40210 19770
rect -40150 19710 -40140 19770
rect -40220 19700 -40140 19710
rect -40180 19650 -40150 19700
rect -40030 19620 -40000 20530
rect -39460 20490 -39430 20540
rect -38940 20490 -38910 20540
rect -39570 20460 -38910 20490
rect -39390 20140 -38690 20180
rect -38500 20170 -38470 22330
rect -38270 22080 -38240 24230
rect -38130 24270 -38050 24280
rect -38130 24210 -38120 24270
rect -38060 24210 -38050 24270
rect -38130 24200 -38050 24210
rect -38080 24150 -38050 24200
rect -37940 24120 -37910 25030
rect -37780 23470 -37750 26920
rect -37370 26300 -37340 26350
rect -36850 26300 -36820 26350
rect -37480 26270 -36820 26300
rect -36410 26000 -36380 28090
rect -36230 27890 -36150 27900
rect -36230 27830 -36220 27890
rect -36160 27830 -36150 27890
rect -36230 27820 -36150 27830
rect -37310 25970 -36600 26000
rect -36410 25990 -36330 26000
rect -37310 25960 -36520 25970
rect -37310 25900 -36590 25960
rect -36530 25900 -36520 25960
rect -37310 25890 -36520 25900
rect -36410 25930 -36400 25990
rect -36340 25930 -36330 25990
rect -36410 25920 -36330 25930
rect -37310 25860 -36600 25890
rect -36600 25620 -36520 25630
rect -36600 25580 -36590 25620
rect -37110 25560 -36590 25580
rect -36530 25560 -36520 25620
rect -37110 25550 -36520 25560
rect -37110 25500 -37080 25550
rect -36600 25500 -36570 25550
rect -37490 24070 -37460 24340
rect -37370 24070 -37340 24120
rect -36850 24070 -36820 24120
rect -37490 24040 -36820 24070
rect -37490 23660 -37460 24040
rect -36410 23760 -36380 25920
rect -36180 25660 -36150 27820
rect -36040 27860 -35960 27870
rect -36040 27800 -36030 27860
rect -35970 27800 -35960 27860
rect -34510 27860 -34430 27870
rect -34510 27820 -34500 27860
rect -36040 27790 -35960 27800
rect -35020 27800 -34500 27820
rect -34440 27800 -34430 27860
rect -35020 27790 -34430 27800
rect -36000 27740 -35970 27790
rect -35690 27780 -35610 27790
rect -35690 27740 -35680 27780
rect -35870 27720 -35680 27740
rect -35620 27720 -35610 27780
rect -35020 27730 -34990 27790
rect -34510 27730 -34480 27790
rect -35870 27710 -35610 27720
rect -35960 25970 -35900 26000
rect -36040 25960 -35900 25970
rect -36040 25900 -36030 25960
rect -35970 25900 -35900 25960
rect -36040 25890 -35900 25900
rect -35960 25860 -35900 25890
rect -36230 25650 -36150 25660
rect -36230 25590 -36220 25650
rect -36160 25590 -36150 25650
rect -36230 25580 -36150 25590
rect -36040 25620 -35960 25630
rect -36040 25560 -36030 25620
rect -35970 25560 -35960 25620
rect -36040 25550 -35960 25560
rect -36000 25500 -35970 25550
rect -35850 25470 -35820 26380
rect -35280 26300 -35250 26350
rect -34760 26300 -34730 26350
rect -35390 26270 -34730 26300
rect -34320 26000 -34290 28090
rect -34140 27890 -34060 27900
rect -34140 27830 -34130 27890
rect -34070 27830 -34060 27890
rect -34140 27820 -34060 27830
rect -35220 25970 -34510 26000
rect -34320 25990 -34210 26000
rect -35220 25960 -34430 25970
rect -35220 25900 -34500 25960
rect -34440 25900 -34430 25960
rect -35220 25890 -34430 25900
rect -34320 25930 -34280 25990
rect -34220 25930 -34210 25990
rect -34320 25920 -34210 25930
rect -35220 25860 -34510 25890
rect -34510 25620 -34430 25630
rect -34510 25580 -34500 25620
rect -35020 25560 -34500 25580
rect -34440 25560 -34430 25620
rect -35020 25550 -34430 25560
rect -35020 25500 -34990 25550
rect -34500 25500 -34470 25550
rect -37310 23730 -35900 23760
rect -35750 23660 -35720 24340
rect -35390 24070 -35360 24340
rect -35280 24070 -35250 24120
rect -34760 24070 -34730 24120
rect -35390 24040 -34730 24070
rect -35390 23660 -35360 24040
rect -34320 23760 -34290 25920
rect -34090 25660 -34060 27820
rect -33950 27860 -33870 27870
rect -33950 27800 -33940 27860
rect -33880 27800 -33870 27860
rect -33950 27790 -33870 27800
rect -33910 27730 -33880 27790
rect -33780 27710 -33570 27740
rect -33870 25970 -33810 26000
rect -33950 25960 -33810 25970
rect -33950 25900 -33940 25960
rect -33880 25900 -33810 25960
rect -33950 25890 -33810 25900
rect -33870 25860 -33810 25890
rect -34140 25650 -34060 25660
rect -34140 25590 -34130 25650
rect -34070 25590 -34060 25650
rect -34140 25580 -34060 25590
rect -33950 25620 -33870 25630
rect -33950 25560 -33940 25620
rect -33880 25560 -33870 25620
rect -33950 25550 -33870 25560
rect -33910 25500 -33880 25550
rect -33760 25470 -33730 26380
rect -35220 23730 -33810 23760
rect -34320 23670 -34060 23700
rect -34320 23660 -34290 23670
rect -37490 23630 -34290 23660
rect -34090 23660 -34060 23670
rect -33660 23660 -33630 24340
rect -34260 23630 -34180 23640
rect -34090 23630 -33630 23660
rect -34260 23590 -34250 23630
rect -37200 23570 -34250 23590
rect -34190 23570 -34180 23630
rect -37200 23560 -34180 23570
rect -33660 23560 -33630 23630
rect -33600 23620 -33570 27710
rect -32140 27120 -32110 28270
rect -32080 27290 -32050 28330
rect -31970 27650 -31870 27680
rect -31760 27650 -31560 27680
rect -31970 27420 -31940 27650
rect -32020 27410 -31940 27420
rect -32020 27350 -32010 27410
rect -31950 27350 -31940 27410
rect -32020 27340 -31940 27350
rect -32080 27260 -31800 27290
rect -31590 27200 -31560 27650
rect -31190 27290 -31160 27680
rect -30470 27290 -30440 27680
rect -31190 27260 -31080 27290
rect -30470 27260 -30360 27290
rect -31590 27190 -31510 27200
rect -31590 27130 -31580 27190
rect -31520 27130 -31510 27190
rect -31590 27120 -31510 27130
rect -32140 27090 -31560 27120
rect -32140 24840 -32110 27090
rect -32140 24830 -31950 24840
rect -32140 24810 -32020 24830
rect -32030 24770 -32020 24810
rect -31960 24770 -31950 24830
rect -32030 24760 -31950 24770
rect -30000 24730 -29600 29560
rect -29540 29550 -29140 29560
rect -29540 29490 -29530 29550
rect -29470 29490 -29140 29550
rect -29540 29270 -29140 29490
rect -29000 29410 -27510 29420
rect -29000 29380 -27580 29410
rect -27590 29350 -27580 29380
rect -27520 29350 -27510 29410
rect -27590 29340 -27510 29350
rect -29540 29070 -27740 29270
rect -29540 25360 -29140 29070
rect -29060 29030 -29020 29070
rect -28810 29030 -28770 29070
rect -28550 29030 -28510 29070
rect -28300 29030 -28260 29070
rect -28040 29030 -28000 29070
rect -27780 29030 -27740 29070
rect -28940 27600 -28900 27640
rect -28680 27600 -28640 27640
rect -28420 27600 -28380 27640
rect -28170 27600 -28130 27640
rect -27910 27600 -27870 27640
rect -27660 27600 -27620 27640
rect -28940 27400 -26680 27600
rect -29000 27260 -27590 27290
rect -29000 27250 -27510 27260
rect -29000 27190 -27580 27250
rect -27520 27190 -27510 27250
rect -29000 27180 -27510 27190
rect -29000 27150 -27590 27180
rect -27080 27040 -26680 27400
rect -28940 26840 -26680 27040
rect -28940 26790 -28900 26840
rect -28680 26790 -28640 26840
rect -28430 26790 -28390 26840
rect -28170 26790 -28130 26840
rect -27910 26790 -27870 26840
rect -27660 26790 -27620 26840
rect -29060 25360 -29020 25410
rect -28810 25360 -28770 25410
rect -28520 25400 -28510 25410
rect -28550 25360 -28510 25400
rect -28300 25400 -28290 25410
rect -28010 25400 -28000 25410
rect -27750 25400 -27740 25410
rect -28300 25360 -28260 25400
rect -28040 25360 -28000 25400
rect -27780 25360 -27740 25400
rect -29540 25160 -27740 25360
rect -27590 25090 -27510 25100
rect -27590 25050 -27580 25090
rect -29000 25030 -27580 25050
rect -27520 25030 -27510 25090
rect -29000 25020 -27510 25030
rect -29000 25010 -27680 25020
rect -32390 24690 -31940 24720
rect -31720 24700 -29600 24730
rect -33600 23590 -33510 23620
rect -37780 23460 -37700 23470
rect -37780 23400 -37770 23460
rect -37710 23400 -37700 23460
rect -37780 23390 -37700 23400
rect -38050 22380 -37990 22410
rect -38130 22370 -37990 22380
rect -38130 22310 -38120 22370
rect -38060 22310 -37990 22370
rect -38130 22300 -37990 22310
rect -38050 22270 -37990 22300
rect -38320 22070 -38240 22080
rect -38320 22010 -38310 22070
rect -38250 22010 -38240 22070
rect -38320 22000 -38240 22010
rect -38500 20160 -38420 20170
rect -39390 20130 -38610 20140
rect -39390 20070 -38680 20130
rect -38620 20070 -38610 20130
rect -39390 20060 -38610 20070
rect -38500 20100 -38490 20160
rect -38430 20100 -38420 20160
rect -38500 20090 -38420 20100
rect -39390 20040 -38690 20060
rect -38690 19800 -38610 19810
rect -38690 19760 -38680 19800
rect -39200 19740 -38680 19760
rect -38620 19740 -38610 19800
rect -39200 19730 -38610 19740
rect -39200 19680 -39170 19730
rect -38690 19680 -38660 19730
rect -40590 17980 -40510 17990
rect -40590 17920 -40580 17980
rect -40520 17920 -40510 17980
rect -40590 17910 -40510 17920
rect -41490 17880 -40080 17910
rect -39940 17840 -39910 19170
rect -39570 18250 -39540 19190
rect -39460 18250 -39430 18300
rect -38940 18250 -38910 18300
rect -39570 18220 -38910 18250
rect -39570 17840 -39540 18220
rect -38500 17940 -38470 20090
rect -38270 19840 -38240 22000
rect -38130 22040 -38050 22050
rect -38130 21980 -38120 22040
rect -38060 21980 -38050 22040
rect -38130 21970 -38050 21980
rect -38080 21920 -38050 21970
rect -37940 21890 -37910 22800
rect -38050 20140 -37990 20180
rect -38130 20130 -37990 20140
rect -38130 20070 -38120 20130
rect -38060 20070 -37990 20130
rect -38130 20060 -37990 20070
rect -38050 20030 -37990 20060
rect -38320 19830 -38240 19840
rect -38320 19770 -38310 19830
rect -38250 19770 -38240 19830
rect -38320 19760 -38240 19770
rect -38130 19800 -38050 19810
rect -38130 19740 -38120 19800
rect -38060 19740 -38050 19800
rect -38130 19730 -38050 19740
rect -38080 19680 -38050 19730
rect -37940 19650 -37910 20560
rect -39400 17910 -37990 17940
rect -37850 17840 -37820 19190
rect -37700 18390 -37620 18400
rect -37700 18330 -37690 18390
rect -37630 18350 -37620 18390
rect -37200 18350 -37170 23560
rect -33660 23530 -33570 23560
rect -33710 23490 -33630 23500
rect -33710 23480 -33700 23490
rect -36990 23450 -33700 23480
rect -36990 23270 -36950 23450
rect -33710 23430 -33700 23450
rect -33640 23430 -33630 23490
rect -33710 23420 -33630 23430
rect -33600 23380 -33570 23530
rect -33660 23350 -33570 23380
rect -34970 23320 -33850 23350
rect -36990 23130 -36960 23270
rect -36120 23230 -36040 23240
rect -36120 23210 -36110 23230
rect -36150 23170 -36110 23210
rect -36050 23170 -36040 23230
rect -36150 23160 -36040 23170
rect -36990 22880 -36950 23130
rect -36110 21780 -36010 21810
rect -36990 21060 -36960 21780
rect -36160 21460 -36130 21490
rect -36160 21450 -36050 21460
rect -36160 21390 -36120 21450
rect -36060 21390 -36050 21450
rect -36160 21380 -36050 21390
rect -36160 21350 -36130 21380
rect -34970 21260 -34940 23320
rect -34870 22200 -34840 22750
rect -34870 21380 -34840 21930
rect -34870 20560 -34840 21110
rect -36010 19990 -35980 20130
rect -36110 19960 -35980 19990
rect -36120 19680 -36040 19690
rect -36150 19630 -36110 19680
rect -36120 19620 -36110 19630
rect -36050 19620 -36040 19680
rect -36120 19610 -36040 19620
rect -36010 19570 -35980 19960
rect -34870 19750 -34840 20300
rect -36170 19540 -34950 19570
rect -36120 19240 -36040 19250
rect -36120 19220 -36110 19240
rect -36150 19180 -36110 19220
rect -36050 19180 -36040 19240
rect -36150 19170 -36040 19180
rect -34870 18930 -34840 19480
rect -37630 18330 -37170 18350
rect -37700 18320 -37170 18330
rect -39940 17810 -39390 17840
rect -38720 17810 -38120 17840
rect -37900 17810 -37820 17840
rect -37770 18250 -37270 18280
rect -41660 17780 -41480 17810
rect -40820 17780 -40210 17810
rect -39990 17780 -39910 17810
rect -41660 17060 -41630 17780
rect -40590 17740 -40510 17750
rect -40590 17680 -40580 17740
rect -40520 17680 -40510 17740
rect -40590 17670 -40510 17680
rect -40590 17340 -40560 17670
rect -37770 17470 -37740 18250
rect -37700 18180 -37620 18190
rect -37700 18120 -37690 18180
rect -37630 18140 -37620 18180
rect -37300 18140 -37270 18250
rect -37630 18120 -37530 18140
rect -37700 18110 -37530 18120
rect -37500 18110 -37270 18140
rect -34870 18110 -34840 18660
rect -37560 17930 -37530 18110
rect -36110 17790 -35980 17820
rect -37390 17470 -37360 17650
rect -36990 17470 -36960 17790
rect -37770 17440 -37440 17470
rect -37390 17440 -36960 17470
rect -36150 17500 -36040 17510
rect -36150 17460 -36110 17500
rect -36120 17440 -36110 17460
rect -36050 17440 -36040 17500
rect -39870 17340 -39390 17370
rect -39230 17340 -38880 17370
rect -38720 17340 -38020 17370
rect -41320 17310 -40120 17340
rect -40080 17310 -39840 17340
rect -40590 17250 -40560 17310
rect -40590 17240 -40510 17250
rect -40590 17180 -40580 17240
rect -40520 17180 -40510 17240
rect -40590 17170 -40510 17180
rect -39870 17140 -39840 17310
rect -38580 17210 -38500 17220
rect -38580 17170 -38570 17210
rect -41290 17110 -40150 17140
rect -41290 16950 -41260 17110
rect -40780 16950 -40750 17110
rect -40590 17070 -40510 17080
rect -40590 17010 -40580 17070
rect -40520 17010 -40510 17070
rect -40590 17000 -40510 17010
rect -41660 15410 -41630 15450
rect -41550 15410 -41520 15570
rect -41030 15410 -41000 15570
rect -41660 15380 -41000 15410
rect -41660 15110 -41630 15380
rect -40590 15210 -40560 17000
rect -40180 16950 -40150 17110
rect -40050 17110 -39840 17140
rect -40050 16950 -40020 17110
rect -39940 15230 -39910 15460
rect -39990 15220 -39910 15230
rect -41520 15180 -40120 15210
rect -39990 15160 -39980 15220
rect -39920 15160 -39910 15220
rect -39990 15150 -39910 15160
rect -39940 15110 -39910 15150
rect -41660 15080 -41480 15110
rect -40810 15080 -40210 15110
rect -39990 15080 -39910 15110
rect -41630 15000 -41600 15080
rect -39870 15070 -39840 17110
rect -39200 17150 -38570 17170
rect -38510 17150 -38500 17210
rect -39200 17140 -38500 17150
rect -39200 16970 -39170 17140
rect -38680 16970 -38650 17140
rect -39570 15440 -39540 15490
rect -39460 15440 -39430 15600
rect -38940 15440 -38910 15600
rect -39570 15410 -38910 15440
rect -39570 15190 -39540 15410
rect -38470 15240 -38440 17340
rect -38210 17210 -38130 17220
rect -38210 17150 -38200 17210
rect -38140 17170 -38130 17210
rect -37770 17170 -37740 17440
rect -36120 17430 -36040 17440
rect -36010 17400 -35980 17680
rect -37350 17370 -36900 17400
rect -36170 17370 -34960 17400
rect -34870 17300 -34840 17830
rect -38140 17150 -38060 17170
rect -38210 17140 -38060 17150
rect -38090 16980 -38060 17140
rect -37960 17140 -37740 17170
rect -37960 16980 -37930 17140
rect -37770 15970 -37740 17140
rect -36120 17070 -36040 17080
rect -36120 17050 -36110 17070
rect -36990 17010 -36910 17040
rect -36150 17010 -36110 17050
rect -36050 17010 -36040 17070
rect -36990 16710 -36960 17010
rect -36150 17000 -36040 17010
rect -37770 15940 -37520 15970
rect -37550 15910 -37470 15940
rect -37550 15720 -37520 15910
rect -39240 15210 -38020 15240
rect -39570 15180 -39490 15190
rect -39570 15120 -39560 15180
rect -39500 15140 -39490 15180
rect -37850 15140 -37820 15490
rect -37550 15330 -37520 15460
rect -37550 15300 -37470 15330
rect -37390 15300 -37360 15480
rect -36990 15300 -36960 15630
rect -36120 15620 -35980 15650
rect -37390 15270 -36890 15300
rect -36010 15230 -35980 15520
rect -34970 15230 -34940 17140
rect -34870 16480 -34840 17020
rect -34870 15660 -34840 16200
rect -37350 15200 -36890 15230
rect -36170 15200 -34940 15230
rect -39500 15120 -39390 15140
rect -39570 15110 -39390 15120
rect -38720 15110 -38120 15140
rect -37900 15110 -37820 15140
rect -34970 15110 -34940 15200
rect -34870 15070 -34840 15380
rect -34780 15180 -34750 23230
rect -33990 17300 -33960 22750
rect -33880 21250 -33850 23320
rect -33660 18780 -33630 23350
rect -33540 20710 -33510 23590
rect -32390 21580 -32360 24690
rect -32090 24590 -31090 24620
rect -30470 24590 -30360 24630
rect -32090 24010 -32060 24590
rect -32030 24330 -31950 24340
rect -32030 24270 -32020 24330
rect -31960 24290 -31950 24330
rect -31960 24270 -31880 24290
rect -32030 24260 -31880 24270
rect -31780 24260 -31570 24290
rect -32090 23980 -31810 24010
rect -31600 23500 -31570 24260
rect -31200 24010 -31170 24590
rect -30470 24340 -30440 24590
rect -31060 24310 -30430 24340
rect -30310 24320 -30280 24700
rect -30000 24560 -29600 24700
rect -27080 24770 -26680 26840
rect -21350 24850 -21240 24870
rect -21350 24780 -21330 24850
rect -21260 24780 -21240 24850
rect -27080 24750 -26570 24770
rect -21350 24760 -21240 24780
rect -21020 24820 -20910 24840
rect -27080 24680 -26660 24750
rect -26590 24680 -26570 24750
rect -21020 24750 -21000 24820
rect -20930 24750 -20910 24820
rect -21020 24730 -20910 24750
rect -27080 24660 -26570 24680
rect -29380 24620 -27120 24630
rect -29380 24600 -27190 24620
rect -27200 24560 -27190 24600
rect -27130 24560 -27120 24620
rect -30000 24390 -27360 24560
rect -27200 24550 -27120 24560
rect -30470 24030 -30440 24310
rect -31200 23980 -31090 24010
rect -30470 23990 -30360 24030
rect -31200 23640 -31170 23980
rect -31200 23630 -31120 23640
rect -31200 23570 -31190 23630
rect -31130 23570 -31120 23630
rect -31200 23560 -31120 23570
rect -31650 23490 -31570 23500
rect -31650 23430 -31640 23490
rect -31580 23430 -31570 23490
rect -31650 23420 -31570 23430
rect -31600 23300 -31570 23420
rect -30000 23510 -29520 24390
rect -29440 24340 -29400 24390
rect -29190 24340 -29150 24390
rect -28930 24340 -28890 24390
rect -28680 24340 -28640 24390
rect -28420 24340 -28380 24390
rect -28160 24340 -28120 24390
rect -27910 24340 -27870 24390
rect -27650 24340 -27610 24390
rect -27400 24340 -27360 24390
rect -29310 24230 -29270 24270
rect -29060 24230 -29020 24270
rect -28800 24230 -28760 24270
rect -28550 24230 -28510 24270
rect -28290 24230 -28250 24270
rect -28030 24230 -27990 24270
rect -27780 24230 -27740 24270
rect -27520 24230 -27480 24270
rect -27270 24230 -27230 24270
rect -27080 24230 -26680 24660
rect -29310 24060 -26680 24230
rect -29380 23990 -27200 24020
rect -29380 23980 -27120 23990
rect -29380 23920 -27190 23980
rect -27130 23920 -27120 23980
rect -29380 23910 -27120 23920
rect -29380 23880 -27200 23910
rect -27080 23840 -26680 24060
rect -29310 23670 -26680 23840
rect -29310 23630 -29270 23670
rect -29060 23630 -29020 23670
rect -28800 23630 -28760 23670
rect -28550 23630 -28510 23670
rect -28290 23630 -28250 23670
rect -28040 23630 -28000 23670
rect -27780 23630 -27740 23670
rect -27520 23630 -27480 23670
rect -27270 23630 -27230 23670
rect -29440 23510 -29400 23560
rect -29190 23510 -29150 23560
rect -28930 23510 -28890 23560
rect -28670 23510 -28630 23560
rect -28420 23510 -28380 23560
rect -28160 23510 -28120 23560
rect -27910 23510 -27870 23560
rect -27650 23510 -27610 23560
rect -27400 23510 -27360 23560
rect -30000 23340 -27360 23510
rect -27200 23340 -27120 23350
rect -27200 23300 -27190 23340
rect -31600 23280 -27190 23300
rect -27130 23280 -27120 23340
rect -31600 23270 -27120 23280
rect -29380 23260 -27290 23270
rect -32390 21570 -28960 21580
rect -32390 21550 -29430 21570
rect -29440 21510 -29430 21550
rect -29370 21550 -28960 21570
rect -28650 21550 -28110 21580
rect -29370 21510 -29360 21550
rect -29440 21500 -29360 21510
rect -28580 21430 -28550 21550
rect -28690 21400 -28550 21430
rect -28210 21430 -28180 21550
rect -28210 21400 -28070 21430
rect -27520 21170 -27490 23260
rect -29270 21140 -28920 21170
rect -27840 21140 -27490 21170
rect -29270 21030 -29240 21140
rect -29270 21000 -28890 21030
rect -28720 21000 -28040 21030
rect -33540 20700 -29300 20710
rect -33540 20680 -29370 20700
rect -29380 20640 -29370 20680
rect -29310 20640 -29300 20700
rect -29380 20630 -29300 20640
rect -33660 18750 -32260 18780
rect -33860 18690 -32330 18720
rect -33990 16910 -33960 17010
rect -33340 16910 -33310 17980
rect -33990 16880 -33310 16910
rect -33990 16480 -33960 16880
rect -33990 15660 -33960 16200
rect -39870 15040 -34840 15070
rect -36190 14900 -36110 14910
rect -36190 14840 -36180 14900
rect -36120 14860 -36110 14900
rect -34780 14860 -34750 15160
rect -36120 14840 -34070 14860
rect -36190 14830 -34070 14840
rect -35110 10720 -35080 11790
rect -35220 10700 -35080 10720
rect -35220 10630 -35200 10700
rect -35130 10630 -35080 10700
rect -35220 10610 -35080 10630
rect -35110 8770 -35080 10610
rect -34100 9750 -34070 14830
rect -33340 10900 -33310 16880
rect -34620 9720 -34070 9750
rect -34620 9590 -34590 9720
rect -34620 9560 -34550 9590
rect -33340 9560 -33260 9590
rect -34620 9350 -34590 9560
rect -33340 9500 -33310 9560
rect -33750 9470 -33310 9500
rect -33750 9350 -33720 9470
rect -33340 9350 -33310 9470
rect -34620 8870 -34590 9070
rect -34620 8840 -34550 8870
rect -33630 8770 -33600 8990
rect -33340 8870 -33310 9070
rect -33340 8840 -33260 8870
rect -33220 8830 -33190 18500
rect -32460 18270 -32430 18660
rect -32460 17450 -32430 17980
rect -32460 16630 -32430 17160
rect -32360 16500 -32330 18690
rect -32290 18030 -32260 18750
rect -29330 18610 -29300 20630
rect -29270 20340 -29240 21000
rect -29030 20510 -28480 20540
rect -29270 20310 -28660 20340
rect -29090 20150 -29060 20310
rect -28690 20150 -28660 20310
rect -28890 18610 -28860 18770
rect -29330 18580 -28860 18610
rect -28510 18410 -28480 20510
rect -28280 20510 -27730 20540
rect -28390 18570 -28310 18580
rect -28390 18510 -28380 18570
rect -28320 18530 -28310 18570
rect -28280 18530 -28250 20510
rect -27520 20340 -27490 21140
rect -28100 20310 -27490 20340
rect -27460 20700 -27380 20710
rect -27460 20640 -27450 20700
rect -27390 20640 -27380 20700
rect -27460 20630 -27380 20640
rect -28100 20150 -28070 20310
rect -27700 20150 -27670 20310
rect -27900 18600 -27870 18760
rect -27460 18600 -27430 20630
rect -27900 18570 -27430 18600
rect -28320 18510 -28250 18530
rect -28390 18500 -28250 18510
rect -28390 18450 -28310 18460
rect -28390 18410 -28380 18450
rect -29030 18390 -28380 18410
rect -28320 18390 -28310 18450
rect -29030 18380 -28310 18390
rect -28280 18410 -28250 18500
rect -28280 18380 -27730 18410
rect -32230 18130 -32150 18140
rect -32230 18070 -32220 18130
rect -32160 18090 -32150 18130
rect -32060 18130 -31980 18140
rect -32060 18090 -32050 18130
rect -32160 18070 -32050 18090
rect -31990 18070 -31980 18130
rect -32230 18060 -31980 18070
rect -28710 18030 -28670 18310
rect -28660 18270 -28050 18310
rect -28500 18230 -28420 18240
rect -28500 18170 -28490 18230
rect -28430 18170 -28420 18230
rect -28500 18160 -28420 18170
rect -28390 18230 -28310 18240
rect -28390 18170 -28380 18230
rect -28320 18170 -28310 18230
rect -28390 18160 -28310 18170
rect -32290 18000 -28670 18030
rect -32170 17950 -32090 17960
rect -32170 17890 -32160 17950
rect -32100 17890 -32090 17950
rect -32170 17880 -32090 17890
rect -32120 17290 -32090 17880
rect -28630 17900 -28550 17910
rect -28630 17860 -28620 17900
rect -30380 17830 -30290 17860
rect -28720 17840 -28620 17860
rect -28560 17860 -28550 17900
rect -28560 17840 -28480 17860
rect -28720 17830 -28480 17840
rect -28630 17400 -28550 17410
rect -28630 17360 -28620 17400
rect -32010 17340 -28620 17360
rect -28560 17340 -28550 17400
rect -32010 17330 -28550 17340
rect -32010 17180 -31970 17330
rect -28690 17180 -28660 17330
rect -32460 15810 -32430 16340
rect -32460 15000 -32430 15530
rect -32460 14170 -32430 14700
rect -32120 14200 -32090 14290
rect -30350 14200 -30320 14400
rect -28620 14240 -28540 14250
rect -28620 14200 -28610 14240
rect -32190 14180 -28610 14200
rect -28550 14180 -28540 14240
rect -32190 14170 -28540 14180
rect -32460 13360 -32430 13890
rect -32190 13350 -32160 14170
rect -30380 13720 -30290 13750
rect -28720 13740 -28550 13750
rect -28720 13720 -28620 13740
rect -28630 13680 -28620 13720
rect -28560 13700 -28550 13740
rect -28510 13700 -28480 17830
rect -28560 13680 -28480 13700
rect -28630 13670 -28480 13680
rect -32190 13340 -28550 13350
rect -32190 13320 -28620 13340
rect -32460 12540 -32430 13070
rect -32460 11720 -32430 12250
rect -32460 10910 -32430 11440
rect -32460 10250 -32430 10620
rect -32350 10250 -32320 12380
rect -32460 10220 -32320 10250
rect -32460 9360 -32430 10220
rect -32350 9520 -32320 10220
rect -32190 9520 -32160 13320
rect -28630 13280 -28620 13320
rect -28560 13280 -28550 13340
rect -28630 13270 -28550 13280
rect -28630 13220 -28550 13230
rect -28630 13180 -28620 13220
rect -30380 13150 -30290 13180
rect -28720 13160 -28620 13180
rect -28560 13180 -28550 13220
rect -28510 13180 -28480 13670
rect -28560 13160 -28480 13180
rect -28720 13150 -28480 13160
rect -28630 12720 -28550 12730
rect -28630 12680 -28620 12720
rect -32010 12660 -28620 12680
rect -28560 12660 -28550 12720
rect -32010 12650 -28550 12660
rect -32010 12500 -31980 12650
rect -28690 12500 -28660 12650
rect -32120 9520 -32090 9610
rect -30350 9520 -30320 9720
rect -28620 9560 -28540 9570
rect -28620 9520 -28610 9560
rect -32350 9500 -28610 9520
rect -28550 9500 -28540 9560
rect -32350 9490 -28540 9500
rect -32350 9430 -32320 9490
rect -28510 9070 -28480 13150
rect -30380 9040 -30290 9070
rect -28720 9060 -28480 9070
rect -28720 9040 -28620 9060
rect -28630 9000 -28620 9040
rect -28560 9040 -28480 9060
rect -28450 17410 -28420 18160
rect -28340 17520 -28310 18160
rect -28090 18030 -28050 18270
rect -28090 18000 -24570 18030
rect -28210 17900 -28130 17910
rect -28210 17840 -28200 17900
rect -28140 17860 -28130 17900
rect -28140 17840 -28040 17860
rect -28210 17830 -28040 17840
rect -26470 17830 -26380 17860
rect -24600 17630 -24570 18000
rect -24600 17600 -24330 17630
rect -24110 17600 -23610 17630
rect -23390 17600 -22890 17630
rect -22670 17600 -22510 17630
rect -28390 17510 -28310 17520
rect -28390 17450 -28380 17510
rect -28320 17450 -28310 17510
rect -28390 17440 -28310 17450
rect -28450 17400 -28370 17410
rect -28450 17340 -28440 17400
rect -28380 17340 -28370 17400
rect -28450 17330 -28370 17340
rect -28450 12730 -28420 17330
rect -28450 12720 -28370 12730
rect -28450 12660 -28440 12720
rect -28380 12660 -28370 12720
rect -28450 12650 -28370 12660
rect -28340 12680 -28310 17440
rect -24480 17500 -24240 17530
rect -23760 17500 -23520 17530
rect -23040 17500 -22800 17530
rect -28210 17400 -28130 17410
rect -28210 17340 -28200 17400
rect -28140 17360 -28130 17400
rect -24480 17360 -24450 17500
rect -28140 17340 -24450 17360
rect -28210 17330 -24450 17340
rect -23990 17370 -23910 17380
rect -23990 17330 -23980 17370
rect -28100 17180 -28070 17330
rect -24780 17180 -24750 17330
rect -24480 15440 -24450 17330
rect -24170 17310 -23980 17330
rect -23920 17310 -23910 17370
rect -24170 17300 -23910 17310
rect -24170 17140 -24140 17300
rect -24300 15600 -24270 15760
rect -24530 15430 -24450 15440
rect -24530 15370 -24520 15430
rect -24460 15370 -24450 15430
rect -24530 15360 -24450 15370
rect -24410 15570 -24270 15600
rect -24410 15160 -24380 15570
rect -24350 15410 -24240 15420
rect -24350 15350 -24340 15410
rect -24280 15350 -24240 15410
rect -24350 15340 -24240 15350
rect -23760 15270 -23730 17500
rect -23270 17370 -23190 17380
rect -23270 17330 -23260 17370
rect -23450 17310 -23260 17330
rect -23200 17310 -23190 17370
rect -23450 17300 -23190 17310
rect -23450 17140 -23420 17300
rect -23580 15600 -23550 15760
rect -23810 15260 -23730 15270
rect -23810 15200 -23800 15260
rect -23740 15200 -23730 15260
rect -23810 15190 -23730 15200
rect -23690 15570 -23550 15600
rect -23690 15160 -23660 15570
rect -23040 15400 -23010 17500
rect -22540 16140 -22510 17600
rect -22540 16100 -22170 16140
rect -21950 16100 -20770 16130
rect -22370 16040 -22130 16050
rect -22370 15980 -22360 16040
rect -22300 16020 -22130 16040
rect -22080 16030 -21800 16060
rect -22300 15980 -22290 16020
rect -22370 15970 -22290 15980
rect -22170 15840 -22130 16020
rect -21980 15860 -21870 15870
rect -21980 15800 -21940 15860
rect -21880 15800 -21870 15860
rect -21980 15790 -21870 15800
rect -22860 15540 -22830 15760
rect -22970 15530 -22830 15540
rect -22970 15470 -22960 15530
rect -22900 15510 -22830 15530
rect -22730 15540 -22700 15760
rect -22620 15580 -22540 15590
rect -22620 15540 -22610 15580
rect -22730 15520 -22610 15540
rect -22550 15520 -22540 15580
rect -22730 15510 -22540 15520
rect -22900 15470 -22890 15510
rect -22970 15460 -22890 15470
rect -21830 15400 -21800 16030
rect -21770 15860 -21690 15870
rect -21770 15800 -21760 15860
rect -21700 15800 -21690 15860
rect -21770 15790 -21690 15800
rect -23480 15370 -23240 15400
rect -23270 15270 -23240 15370
rect -23040 15370 -22080 15400
rect -22040 15370 -21800 15400
rect -23270 15260 -23190 15270
rect -23270 15200 -23260 15260
rect -23200 15200 -23190 15260
rect -23270 15190 -23190 15200
rect -23040 15160 -23010 15370
rect -24410 15130 -23010 15160
rect -22970 15200 -22890 15210
rect -22970 15140 -22960 15200
rect -22900 15160 -22890 15200
rect -22900 15140 -20950 15160
rect -22970 15130 -20950 15140
rect -24410 14410 -24380 15130
rect -20980 15000 -20950 15130
rect -22670 14960 -22580 14990
rect -21010 14950 -20950 15000
rect -20980 14400 -20950 14950
rect -28210 14250 -28180 14290
rect -28220 14240 -28140 14250
rect -28220 14180 -28210 14240
rect -28150 14200 -28140 14240
rect -26440 14200 -26410 14400
rect -24300 14370 -20950 14400
rect -24300 14310 -24270 14370
rect -20980 14310 -20950 14370
rect -28150 14180 -26410 14200
rect -28220 14170 -26410 14180
rect -28210 13740 -28040 13750
rect -28210 13680 -28200 13740
rect -28140 13720 -28040 13740
rect -26470 13720 -26380 13750
rect -28140 13680 -28130 13720
rect -28210 13670 -28130 13680
rect -28210 13340 -24380 13350
rect -28210 13280 -28200 13340
rect -28140 13320 -24380 13340
rect -28140 13280 -28130 13320
rect -28210 13270 -28130 13280
rect -28210 13220 -28130 13230
rect -28210 13160 -28200 13220
rect -28140 13180 -28130 13220
rect -28140 13160 -28040 13180
rect -28210 13150 -28040 13160
rect -26470 13150 -26380 13180
rect -24600 12720 -24520 12730
rect -24600 12680 -24590 12720
rect -28340 12660 -24590 12680
rect -24530 12660 -24520 12720
rect -28340 12650 -24520 12660
rect -28560 9000 -28550 9040
rect -28630 8990 -28550 9000
rect -32360 8770 -32330 8990
rect -35110 8740 -34430 8770
rect -33900 8740 -33150 8770
rect -32620 8740 -32330 8770
rect -35260 8710 -35180 8720
rect -35260 8650 -35250 8710
rect -35190 8650 -35180 8710
rect -35260 8640 -35180 8650
rect -35210 4870 -35180 8640
rect -28620 8600 -28540 8610
rect -29560 8570 -28610 8600
rect -28620 8540 -28610 8570
rect -28550 8540 -28540 8600
rect -28620 8530 -28540 8540
rect -34960 8470 -28480 8500
rect -28630 8040 -28550 8050
rect -28630 8000 -28620 8040
rect -35030 7980 -28620 8000
rect -28560 7980 -28550 8040
rect -35030 7970 -28550 7980
rect -35030 7810 -35000 7970
rect -34630 7810 -34600 7970
rect -34240 7810 -34210 7970
rect -33840 7810 -33810 7970
rect -33440 7810 -33410 7970
rect -33050 7810 -33020 7970
rect -32650 7810 -32620 7970
rect -32260 7810 -32230 7970
rect -31860 7810 -31830 7970
rect -31460 7810 -31430 7970
rect -31070 7810 -31040 7970
rect -30670 7810 -30640 7970
rect -30280 7810 -30250 7970
rect -29880 7810 -29850 7970
rect -29480 7810 -29450 7970
rect -29090 7810 -29060 7970
rect -28690 7810 -28660 7970
rect -34830 4870 -34800 5030
rect -34430 4870 -34400 5030
rect -34040 4870 -34010 5030
rect -33640 4870 -33610 5030
rect -33250 4870 -33220 5030
rect -32850 4870 -32820 5030
rect -32450 4870 -32420 5030
rect -32060 4870 -32030 5030
rect -31660 4870 -31630 5030
rect -31270 4870 -31240 5030
rect -30870 4870 -30840 5030
rect -30480 4870 -30450 5030
rect -30080 4870 -30050 5030
rect -29680 4870 -29650 5030
rect -29290 4870 -29260 5030
rect -28890 4870 -28860 5030
rect -35210 4860 -28540 4870
rect -35210 4840 -28610 4860
rect -35210 170 -35180 4840
rect -28620 4800 -28610 4840
rect -28550 4800 -28540 4860
rect -28620 4790 -28540 4800
rect -28510 4370 -28480 8470
rect -34970 4360 -28480 4370
rect -34970 4340 -28550 4360
rect -28560 4300 -28550 4340
rect -28490 4300 -28480 4360
rect -28560 4290 -28480 4300
rect -28510 4110 -28480 4290
rect -28560 4100 -28480 4110
rect -35150 4030 -35040 4050
rect -28560 4040 -28550 4100
rect -28490 4040 -28480 4100
rect -28560 4030 -28480 4040
rect -28450 8050 -28420 12650
rect -28340 8160 -28310 12650
rect -28100 12500 -28070 12650
rect -24780 12500 -24750 12650
rect -22640 11450 -22610 11530
rect -24410 11420 -22610 11450
rect -20980 10890 -20950 11530
rect -24600 10850 -24240 10880
rect -22670 10850 -22580 10880
rect -21010 10850 -20950 10890
rect -28210 9570 -28180 9610
rect -28220 9560 -28140 9570
rect -28220 9500 -28210 9560
rect -28150 9520 -28140 9560
rect -26440 9520 -26410 9720
rect -28150 9500 -26410 9520
rect -28220 9490 -26410 9500
rect -24600 9070 -24570 10850
rect -20800 10580 -20770 16100
rect -28210 9060 -28040 9070
rect -28210 9000 -28200 9060
rect -28140 9040 -28040 9060
rect -26470 9040 -26380 9070
rect -24810 9040 -24570 9070
rect -21650 10550 -20770 10580
rect -28140 9000 -28130 9040
rect -28210 8990 -28130 9000
rect -28220 8600 -27200 8610
rect -21650 8600 -21620 10550
rect -28220 8540 -28210 8600
rect -28150 8580 -27200 8600
rect -28150 8540 -28140 8580
rect -22630 8570 -21620 8600
rect -28220 8530 -28140 8540
rect -28390 8150 -28310 8160
rect -28390 8090 -28380 8150
rect -28320 8090 -28310 8150
rect -28390 8080 -28310 8090
rect -28450 8040 -28370 8050
rect -28450 7980 -28440 8040
rect -28380 7980 -28370 8040
rect -28450 7970 -28370 7980
rect -35150 3960 -35130 4030
rect -35060 3960 -35040 4030
rect -35150 3940 -35040 3960
rect -35150 3300 -35120 3940
rect -28560 3840 -28480 3850
rect -28560 3800 -28550 3840
rect -34970 3780 -28550 3800
rect -28490 3780 -28480 3840
rect -34970 3770 -28480 3780
rect -28630 3340 -28550 3350
rect -28630 3300 -28620 3340
rect -35150 3280 -28620 3300
rect -28560 3280 -28550 3340
rect -35150 3270 -28550 3280
rect -35030 3110 -35000 3270
rect -34630 3110 -34600 3270
rect -34240 3110 -34210 3270
rect -33840 3110 -33810 3270
rect -33440 3110 -33410 3270
rect -33050 3110 -33020 3270
rect -32650 3110 -32620 3270
rect -32260 3110 -32230 3270
rect -31860 3110 -31830 3270
rect -31460 3110 -31430 3270
rect -31070 3110 -31040 3270
rect -30670 3110 -30640 3270
rect -30280 3110 -30250 3270
rect -29880 3110 -29850 3270
rect -29480 3110 -29450 3270
rect -29090 3110 -29060 3270
rect -28690 3110 -28660 3270
rect -34830 170 -34800 330
rect -34430 170 -34400 330
rect -34040 170 -34010 330
rect -33640 170 -33610 330
rect -33250 170 -33220 330
rect -32850 170 -32820 330
rect -32450 170 -32420 330
rect -32060 170 -32030 330
rect -31660 170 -31630 330
rect -31270 170 -31240 330
rect -30870 170 -30840 330
rect -30480 170 -30450 330
rect -30080 170 -30050 330
rect -29680 170 -29650 330
rect -29290 170 -29260 330
rect -28890 170 -28860 330
rect -35210 160 -28540 170
rect -35210 140 -28610 160
rect -28620 100 -28610 140
rect -28550 100 -28540 160
rect -28620 90 -28540 100
rect -28510 -330 -28480 3770
rect -28450 3350 -28420 7970
rect -28340 3460 -28310 8080
rect -28280 8470 -21790 8500
rect -28280 4370 -28250 8470
rect -28210 8040 -28130 8050
rect -28210 7980 -28200 8040
rect -28140 8000 -28130 8040
rect -28140 7980 -21730 8000
rect -28210 7970 -21730 7980
rect -28100 7810 -28070 7970
rect -27700 7810 -27670 7970
rect -27310 7810 -27280 7970
rect -26910 7810 -26880 7970
rect -26510 7810 -26480 7970
rect -26120 7810 -26090 7970
rect -25720 7810 -25690 7970
rect -25330 7810 -25300 7970
rect -24930 7810 -24900 7970
rect -24530 7810 -24500 7970
rect -24140 7810 -24110 7970
rect -23740 7810 -23710 7970
rect -23350 7810 -23320 7970
rect -22950 7810 -22920 7970
rect -22550 7810 -22520 7970
rect -22160 7810 -22130 7970
rect -21760 7810 -21730 7970
rect -21650 7920 -21620 8570
rect -27900 4870 -27870 5030
rect -27500 4870 -27470 5030
rect -27110 4870 -27080 5030
rect -26710 4870 -26680 5030
rect -26320 4870 -26290 5030
rect -25920 4870 -25890 5030
rect -25520 4870 -25490 5030
rect -25130 4870 -25100 5030
rect -24730 4870 -24700 5030
rect -24340 4870 -24310 5030
rect -23940 4870 -23910 5030
rect -23550 4870 -23520 5030
rect -23150 4870 -23120 5030
rect -22750 4870 -22720 5030
rect -22360 4870 -22330 5030
rect -21960 4870 -21930 5030
rect -28220 4860 -21930 4870
rect -28220 4800 -28210 4860
rect -28150 4840 -21930 4860
rect -28150 4800 -28140 4840
rect -28220 4790 -28140 4800
rect -28280 4360 -21790 4370
rect -28280 4300 -28270 4360
rect -28210 4340 -21790 4360
rect -28210 4300 -28200 4340
rect -28280 4290 -28200 4300
rect -21650 4270 -21620 4920
rect -22630 4240 -21620 4270
rect -21650 3900 -21620 4240
rect -22630 3870 -21620 3900
rect -28390 3450 -28310 3460
rect -28390 3390 -28380 3450
rect -28320 3390 -28310 3450
rect -28390 3380 -28310 3390
rect -28280 3840 -28200 3850
rect -28280 3780 -28270 3840
rect -28210 3800 -28200 3840
rect -28210 3780 -21790 3800
rect -28280 3770 -21790 3780
rect -28450 3340 -28370 3350
rect -28450 3280 -28440 3340
rect -28380 3280 -28370 3340
rect -28450 3270 -28370 3280
rect -34970 -360 -28480 -330
rect -28620 -400 -28540 -390
rect -28620 -430 -28610 -400
rect -29560 -460 -28610 -430
rect -28550 -460 -28540 -400
rect -28620 -470 -28540 -460
rect -28510 -580 -28480 -360
rect -28280 -330 -28250 3770
rect -21650 3520 -21620 3870
rect -21700 3510 -21620 3520
rect -21700 3450 -21690 3510
rect -21630 3450 -21620 3510
rect -21700 3440 -21620 3450
rect -21760 3380 -21550 3410
rect -28210 3340 -28130 3350
rect -28210 3280 -28200 3340
rect -28140 3300 -28130 3340
rect -21760 3300 -21730 3380
rect -28140 3280 -21730 3300
rect -28210 3270 -21730 3280
rect -21700 3340 -21620 3350
rect -21700 3280 -21690 3340
rect -21630 3280 -21620 3340
rect -21700 3270 -21620 3280
rect -28100 3110 -28070 3270
rect -27700 3110 -27670 3270
rect -27310 3110 -27280 3270
rect -26910 3110 -26880 3270
rect -26510 3110 -26480 3270
rect -26120 3110 -26090 3270
rect -25720 3110 -25690 3270
rect -25330 3110 -25300 3270
rect -24930 3110 -24900 3270
rect -24530 3110 -24500 3270
rect -24140 3110 -24110 3270
rect -23740 3110 -23710 3270
rect -23350 3110 -23320 3270
rect -22950 3110 -22920 3270
rect -22550 3110 -22520 3270
rect -22160 3110 -22130 3270
rect -21760 3110 -21730 3270
rect -21650 3220 -21620 3270
rect -27900 170 -27870 330
rect -27500 170 -27470 330
rect -27110 170 -27080 330
rect -26710 170 -26680 330
rect -26320 170 -26290 330
rect -25920 170 -25890 330
rect -25520 170 -25490 330
rect -25130 170 -25100 330
rect -24730 170 -24700 330
rect -24340 170 -24310 330
rect -23940 170 -23910 330
rect -23550 170 -23520 330
rect -23150 170 -23120 330
rect -22750 170 -22720 330
rect -22360 170 -22330 330
rect -21960 170 -21930 330
rect -28220 160 -21930 170
rect -28220 100 -28210 160
rect -28150 140 -21930 160
rect -28150 100 -28140 140
rect -28220 90 -28140 100
rect -28280 -360 -21790 -330
rect -28280 -550 -28250 -360
rect -28220 -400 -28140 -390
rect -28220 -460 -28210 -400
rect -28150 -440 -28140 -400
rect -21650 -430 -21620 210
rect -28150 -460 -27200 -440
rect -22630 -460 -21620 -430
rect -28220 -470 -27200 -460
rect -28310 -580 -28250 -550
rect -28590 -600 -28480 -580
rect -28590 -670 -28570 -600
rect -28500 -670 -28480 -600
rect -28590 -690 -28480 -670
rect -28390 -600 -28280 -580
rect -28390 -670 -28370 -600
rect -28300 -670 -28280 -600
rect -28390 -690 -28280 -670
rect -21580 -760 -21550 3380
rect -15000 -730 -14890 -710
rect -15000 -760 -14980 -730
rect -21580 -790 -14980 -760
rect -15000 -800 -14980 -790
rect -14910 -800 -14890 -730
rect -15000 -820 -14890 -800
<< via1 >>
rect -30140 29490 -30080 29550
rect -40580 29420 -40520 29480
rect -37650 29220 -37590 29280
rect -37420 29220 -37360 29280
rect -32320 28340 -32260 28400
rect -32140 28340 -32080 28400
rect -35680 28200 -35620 28260
rect -36590 27800 -36530 27860
rect -40580 27290 -40520 27350
rect -40580 26730 -40520 26790
rect -40770 26420 -40710 26480
rect -39970 26680 -39910 26740
rect -40520 26390 -40460 26450
rect -40210 26420 -40150 26480
rect -40770 24520 -40710 24580
rect -40580 24550 -40520 24610
rect -40770 24180 -40710 24240
rect -39680 26710 -39620 26770
rect -38680 26450 -38620 26510
rect -40210 24520 -40150 24580
rect -40470 24210 -40410 24270
rect -40770 22290 -40710 22350
rect -40580 22320 -40520 22380
rect -40770 21960 -40710 22020
rect -40210 24180 -40150 24240
rect -38310 26480 -38250 26540
rect -38680 24550 -38620 24610
rect -38490 24580 -38430 24640
rect -38680 24210 -38620 24270
rect -40210 22290 -40150 22350
rect -40470 21990 -40410 22050
rect -40770 20050 -40710 20110
rect -40580 20080 -40520 20140
rect -40770 19710 -40710 19770
rect -40210 21960 -40150 22020
rect -38120 26450 -38060 26510
rect -37880 25550 -37820 25610
rect -38120 24550 -38060 24610
rect -38310 24240 -38250 24300
rect -38680 22310 -38620 22370
rect -38490 22340 -38430 22400
rect -38680 21980 -38620 22040
rect -40210 20050 -40150 20110
rect -40470 19740 -40410 19800
rect -40210 19710 -40150 19770
rect -38120 24210 -38060 24270
rect -36220 27830 -36160 27890
rect -36590 25900 -36530 25960
rect -36400 25930 -36340 25990
rect -36590 25560 -36530 25620
rect -36030 27800 -35970 27860
rect -34500 27800 -34440 27860
rect -35680 27720 -35620 27780
rect -36030 25900 -35970 25960
rect -36220 25590 -36160 25650
rect -36030 25560 -35970 25620
rect -34130 27830 -34070 27890
rect -34500 25900 -34440 25960
rect -34280 25930 -34220 25990
rect -34500 25560 -34440 25620
rect -33940 27800 -33880 27860
rect -33940 25900 -33880 25960
rect -34130 25590 -34070 25650
rect -33940 25560 -33880 25620
rect -34250 23570 -34190 23630
rect -32010 27350 -31950 27410
rect -31580 27130 -31520 27190
rect -32020 24770 -31960 24830
rect -29530 29490 -29470 29550
rect -27580 29350 -27520 29410
rect -27580 27190 -27520 27250
rect -27580 25030 -27520 25090
rect -37770 23400 -37710 23460
rect -38120 22310 -38060 22370
rect -38310 22010 -38250 22070
rect -38680 20070 -38620 20130
rect -38490 20100 -38430 20160
rect -38680 19740 -38620 19800
rect -40580 17920 -40520 17980
rect -38120 21980 -38060 22040
rect -38120 20070 -38060 20130
rect -38310 19770 -38250 19830
rect -38120 19740 -38060 19800
rect -37690 18330 -37630 18390
rect -33700 23430 -33640 23490
rect -36110 23170 -36050 23230
rect -36120 21390 -36060 21450
rect -36110 19620 -36050 19680
rect -36110 19180 -36050 19240
rect -40580 17680 -40520 17740
rect -37690 18120 -37630 18180
rect -36110 17440 -36050 17500
rect -40580 17180 -40520 17240
rect -40580 17010 -40520 17070
rect -39980 15160 -39920 15220
rect -38570 17150 -38510 17210
rect -38200 17150 -38140 17210
rect -36110 17010 -36050 17070
rect -39560 15120 -39500 15180
rect -32020 24270 -31960 24330
rect -21330 24780 -21260 24850
rect -26660 24680 -26590 24750
rect -21000 24750 -20930 24820
rect -27190 24560 -27130 24620
rect -31190 23570 -31130 23630
rect -31640 23430 -31580 23490
rect -27190 23920 -27130 23980
rect -27190 23280 -27130 23340
rect -29430 21510 -29370 21570
rect -29370 20640 -29310 20700
rect -36180 14840 -36120 14900
rect -35200 10630 -35130 10700
rect -28380 18510 -28320 18570
rect -27450 20640 -27390 20700
rect -28380 18390 -28320 18450
rect -32220 18070 -32160 18130
rect -32050 18070 -31990 18130
rect -28490 18170 -28430 18230
rect -28380 18170 -28320 18230
rect -32160 17890 -32100 17950
rect -28620 17840 -28560 17900
rect -28620 17340 -28560 17400
rect -28610 14180 -28550 14240
rect -28620 13680 -28560 13740
rect -28620 13280 -28560 13340
rect -28620 13160 -28560 13220
rect -28620 12660 -28560 12720
rect -28610 9500 -28550 9560
rect -28620 9000 -28560 9060
rect -28200 17840 -28140 17900
rect -28380 17450 -28320 17510
rect -28440 17340 -28380 17400
rect -28440 12660 -28380 12720
rect -28200 17340 -28140 17400
rect -23980 17310 -23920 17370
rect -24520 15370 -24460 15430
rect -24340 15350 -24280 15410
rect -23260 17310 -23200 17370
rect -23800 15200 -23740 15260
rect -22360 15980 -22300 16040
rect -21940 15800 -21880 15860
rect -22960 15470 -22900 15530
rect -22610 15520 -22550 15580
rect -21760 15800 -21700 15860
rect -23260 15200 -23200 15260
rect -22960 15140 -22900 15200
rect -28210 14180 -28150 14240
rect -28200 13680 -28140 13740
rect -28200 13280 -28140 13340
rect -28200 13160 -28140 13220
rect -24590 12660 -24530 12720
rect -35250 8650 -35190 8710
rect -28610 8540 -28550 8600
rect -28620 7980 -28560 8040
rect -28610 4800 -28550 4860
rect -28550 4300 -28490 4360
rect -28550 4040 -28490 4100
rect -28210 9500 -28150 9560
rect -28200 9000 -28140 9060
rect -28210 8540 -28150 8600
rect -28380 8090 -28320 8150
rect -28440 7980 -28380 8040
rect -35130 3960 -35060 4030
rect -28550 3780 -28490 3840
rect -28620 3280 -28560 3340
rect -28610 100 -28550 160
rect -28200 7980 -28140 8040
rect -28210 4800 -28150 4860
rect -28270 4300 -28210 4360
rect -28380 3390 -28320 3450
rect -28270 3780 -28210 3840
rect -28440 3280 -28380 3340
rect -28610 -460 -28550 -400
rect -21690 3450 -21630 3510
rect -28200 3280 -28140 3340
rect -21690 3280 -21630 3340
rect -28210 100 -28150 160
rect -28210 -460 -28150 -400
rect -28570 -670 -28500 -600
rect -28370 -670 -28300 -600
rect -14980 -800 -14910 -730
<< metal2 >>
rect -30150 29550 -30070 29560
rect -30150 29490 -30140 29550
rect -30080 29510 -30070 29550
rect -29540 29550 -29460 29560
rect -29540 29510 -29530 29550
rect -30080 29490 -29530 29510
rect -29470 29490 -29460 29550
rect -40590 29480 -40510 29490
rect -30150 29480 -29460 29490
rect -40590 29420 -40580 29480
rect -40520 29420 -40510 29480
rect -40590 29410 -40510 29420
rect -27590 29410 -27510 29420
rect -40590 27360 -40560 29410
rect -27590 29350 -27580 29410
rect -27520 29350 -27510 29410
rect -27590 29340 -27510 29350
rect -37660 29280 -37580 29290
rect -37660 29220 -37650 29280
rect -37590 29240 -37580 29280
rect -37430 29280 -37350 29290
rect -37430 29240 -37420 29280
rect -37590 29220 -37420 29240
rect -37360 29240 -37350 29280
rect -37360 29220 -32180 29240
rect -37660 29210 -32180 29220
rect -32330 28400 -32250 28410
rect -32330 28340 -32320 28400
rect -32260 28340 -32250 28400
rect -32330 28330 -32250 28340
rect -35690 28260 -35610 28270
rect -35690 28200 -35680 28260
rect -35620 28200 -35610 28260
rect -35690 28190 -35610 28200
rect -36230 27890 -36150 27900
rect -36600 27860 -36520 27870
rect -36600 27800 -36590 27860
rect -36530 27820 -36520 27860
rect -36230 27830 -36220 27890
rect -36160 27830 -36150 27890
rect -36230 27820 -36150 27830
rect -36040 27860 -35960 27870
rect -36040 27820 -36030 27860
rect -36530 27800 -36030 27820
rect -35970 27800 -35960 27860
rect -36600 27790 -35960 27800
rect -35690 27790 -35660 28190
rect -34140 27890 -34060 27900
rect -34510 27860 -34430 27870
rect -34510 27800 -34500 27860
rect -34440 27820 -34430 27860
rect -34140 27830 -34130 27890
rect -34070 27830 -34060 27890
rect -34140 27820 -34060 27830
rect -33950 27860 -33870 27870
rect -33950 27820 -33940 27860
rect -34440 27800 -33940 27820
rect -33880 27800 -33870 27860
rect -34510 27790 -33870 27800
rect -35690 27780 -35610 27790
rect -35690 27720 -35680 27780
rect -35620 27720 -35610 27780
rect -35690 27710 -35610 27720
rect -40590 27350 -40510 27360
rect -40590 27290 -40580 27350
rect -40520 27290 -40510 27350
rect -40590 27280 -40510 27290
rect -40590 26800 -40560 27280
rect -40590 26790 -40510 26800
rect -40590 26730 -40580 26790
rect -40520 26730 -40510 26790
rect -39690 26770 -39610 26780
rect -39690 26750 -39680 26770
rect -40590 26720 -40510 26730
rect -39980 26740 -39680 26750
rect -39980 26680 -39970 26740
rect -39910 26710 -39680 26740
rect -39620 26710 -39610 26770
rect -39910 26700 -39610 26710
rect -39910 26680 -39900 26700
rect -39980 26670 -39900 26680
rect -38320 26540 -38240 26550
rect -38690 26510 -38610 26520
rect -40780 26480 -40140 26490
rect -40780 26420 -40770 26480
rect -40710 26460 -40210 26480
rect -40710 26420 -40700 26460
rect -40780 26410 -40700 26420
rect -40530 26450 -40450 26460
rect -40530 26390 -40520 26450
rect -40460 26390 -40450 26450
rect -40220 26420 -40210 26460
rect -40150 26420 -40140 26480
rect -38690 26450 -38680 26510
rect -38620 26470 -38610 26510
rect -38320 26480 -38310 26540
rect -38250 26480 -38240 26540
rect -38320 26470 -38240 26480
rect -38130 26510 -38050 26520
rect -38130 26470 -38120 26510
rect -38620 26450 -38120 26470
rect -38060 26450 -38050 26510
rect -38690 26440 -38050 26450
rect -40220 26410 -40140 26420
rect -40530 26380 -40450 26390
rect -36410 25990 -36330 26000
rect -36600 25960 -36520 25970
rect -36600 25900 -36590 25960
rect -36530 25920 -36520 25960
rect -36410 25930 -36400 25990
rect -36340 25930 -36330 25990
rect -34290 25990 -34210 26000
rect -36410 25920 -36330 25930
rect -36040 25960 -35960 25970
rect -36040 25920 -36030 25960
rect -36530 25900 -36030 25920
rect -35970 25900 -35960 25960
rect -36600 25890 -35960 25900
rect -34510 25960 -34430 25970
rect -34510 25900 -34500 25960
rect -34440 25920 -34430 25960
rect -34290 25930 -34280 25990
rect -34220 25930 -34210 25990
rect -34290 25920 -34210 25930
rect -33950 25960 -33870 25970
rect -33950 25920 -33940 25960
rect -34440 25900 -33940 25920
rect -33880 25900 -33870 25960
rect -34510 25890 -33870 25900
rect -36230 25650 -36150 25660
rect -36600 25620 -36520 25630
rect -37890 25610 -37810 25620
rect -37890 25550 -37880 25610
rect -37820 25570 -37810 25610
rect -37820 25550 -37680 25570
rect -36600 25560 -36590 25620
rect -36530 25580 -36520 25620
rect -36230 25590 -36220 25650
rect -36160 25590 -36150 25650
rect -34140 25650 -34060 25660
rect -36230 25580 -36150 25590
rect -36040 25620 -35960 25630
rect -36040 25580 -36030 25620
rect -36530 25560 -36030 25580
rect -35970 25560 -35960 25620
rect -36600 25550 -35960 25560
rect -34510 25620 -34430 25630
rect -34510 25560 -34500 25620
rect -34440 25580 -34430 25620
rect -34140 25590 -34130 25650
rect -34070 25590 -34060 25650
rect -34140 25580 -34060 25590
rect -33950 25620 -33870 25630
rect -33950 25580 -33940 25620
rect -34440 25560 -33940 25580
rect -33880 25560 -33870 25620
rect -34510 25550 -33870 25560
rect -37890 25540 -37680 25550
rect -38500 24640 -38420 24650
rect -40590 24610 -40510 24620
rect -40780 24580 -40700 24590
rect -40780 24520 -40770 24580
rect -40710 24540 -40700 24580
rect -40590 24550 -40580 24610
rect -40520 24550 -40510 24610
rect -38690 24610 -38610 24620
rect -40590 24540 -40510 24550
rect -40220 24580 -40140 24590
rect -40220 24540 -40210 24580
rect -40710 24520 -40210 24540
rect -40150 24520 -40140 24580
rect -38690 24550 -38680 24610
rect -38620 24570 -38610 24610
rect -38500 24580 -38490 24640
rect -38430 24580 -38420 24640
rect -38500 24570 -38420 24580
rect -38130 24610 -38050 24620
rect -38130 24570 -38120 24610
rect -38620 24550 -38120 24570
rect -38060 24550 -38050 24610
rect -38690 24540 -38050 24550
rect -40780 24510 -40140 24520
rect -38320 24300 -38240 24310
rect -40480 24270 -40400 24280
rect -40780 24240 -40700 24250
rect -40780 24180 -40770 24240
rect -40710 24200 -40700 24240
rect -40480 24210 -40470 24270
rect -40410 24210 -40400 24270
rect -38690 24270 -38610 24280
rect -40480 24200 -40400 24210
rect -40220 24240 -40140 24250
rect -40220 24200 -40210 24240
rect -40710 24180 -40210 24200
rect -40150 24180 -40140 24240
rect -38690 24210 -38680 24270
rect -38620 24230 -38610 24270
rect -38320 24240 -38310 24300
rect -38250 24240 -38240 24300
rect -38320 24230 -38240 24240
rect -38130 24270 -38050 24280
rect -38130 24230 -38120 24270
rect -38620 24210 -38120 24230
rect -38060 24210 -38050 24270
rect -38690 24200 -38050 24210
rect -40780 24170 -40140 24180
rect -37710 23530 -37680 25540
rect -34260 23630 -34180 23640
rect -34260 23570 -34250 23630
rect -34190 23590 -34180 23630
rect -32330 23590 -32300 28330
rect -34190 23570 -32300 23590
rect -34260 23560 -32300 23570
rect -32210 23590 -32180 29210
rect -32150 28400 -32070 28410
rect -32150 28340 -32140 28400
rect -32080 28340 -32070 28400
rect -32150 28330 -32070 28340
rect -32020 27410 -31940 27420
rect -32020 27350 -32010 27410
rect -31950 27350 -31940 27410
rect -32020 27340 -31940 27350
rect -31970 27060 -31940 27340
rect -27540 27260 -27510 29340
rect -27590 27250 -27510 27260
rect -31590 27190 -31510 27200
rect -31590 27130 -31580 27190
rect -31520 27130 -31510 27190
rect -27590 27190 -27580 27250
rect -27520 27190 -27510 27250
rect -27590 27180 -27510 27190
rect -31590 27120 -31510 27130
rect -31590 27090 -30060 27120
rect -31970 27030 -30120 27060
rect -32030 24830 -31950 24840
rect -32030 24770 -32020 24830
rect -31960 24770 -31950 24830
rect -30150 24800 -30120 27030
rect -30090 24880 -30060 27090
rect -27540 25250 -27510 27180
rect -27540 25220 -21320 25250
rect -27540 25100 -27510 25220
rect -27590 25090 -27510 25100
rect -27590 25030 -27580 25090
rect -27520 25030 -27510 25090
rect -27590 25020 -27510 25030
rect -27540 24880 -27510 25020
rect -30090 24850 -27510 24880
rect -26510 24960 -21380 24990
rect -30150 24770 -27120 24800
rect -32030 24760 -31950 24770
rect -32030 24340 -32000 24760
rect -27150 24630 -27120 24770
rect -26680 24750 -26570 24770
rect -26680 24680 -26660 24750
rect -26590 24680 -26570 24750
rect -26680 24660 -26570 24680
rect -26510 24630 -26480 24960
rect -21410 24730 -21380 24960
rect -21350 24870 -21320 25220
rect -21350 24850 -21240 24870
rect -21350 24780 -21330 24850
rect -21260 24780 -21240 24850
rect -21350 24760 -21240 24780
rect -21020 24820 -20910 24840
rect -21020 24750 -21000 24820
rect -20930 24750 -20910 24820
rect -21020 24730 -20910 24750
rect -21410 24700 -20990 24730
rect -27200 24620 -26480 24630
rect -27200 24560 -27190 24620
rect -27130 24600 -26480 24620
rect -27130 24560 -27120 24600
rect -27200 24550 -27120 24560
rect -32030 24330 -31950 24340
rect -32030 24270 -32020 24330
rect -31960 24270 -31950 24330
rect -32030 24260 -31950 24270
rect -27150 23990 -27120 24550
rect -27200 23980 -27120 23990
rect -27200 23920 -27190 23980
rect -27130 23920 -27120 23980
rect -27200 23910 -27120 23920
rect -31200 23630 -31120 23640
rect -31200 23590 -31190 23630
rect -32210 23570 -31190 23590
rect -31130 23570 -31120 23630
rect -32210 23560 -31120 23570
rect -37710 23500 -33740 23530
rect -37780 23460 -37700 23470
rect -37780 23400 -37770 23460
rect -37710 23420 -37700 23460
rect -37710 23400 -33800 23420
rect -37780 23390 -33800 23400
rect -33830 23290 -33800 23390
rect -33770 23350 -33740 23500
rect -33710 23490 -31570 23500
rect -33710 23430 -33700 23490
rect -33640 23470 -31640 23490
rect -33640 23430 -33630 23470
rect -33710 23420 -33630 23430
rect -31650 23430 -31640 23470
rect -31580 23430 -31570 23490
rect -31650 23420 -31570 23430
rect -27150 23350 -27120 23910
rect -33770 23320 -33570 23350
rect -33830 23260 -33780 23290
rect -36120 23230 -35910 23240
rect -36120 23170 -36110 23230
rect -36050 23210 -35910 23230
rect -36050 23170 -36040 23210
rect -36120 23160 -36040 23170
rect -38500 22400 -38420 22410
rect -40590 22380 -40510 22390
rect -40780 22350 -40700 22360
rect -40780 22290 -40770 22350
rect -40710 22310 -40700 22350
rect -40590 22320 -40580 22380
rect -40520 22320 -40510 22380
rect -38690 22370 -38610 22380
rect -40590 22310 -40510 22320
rect -40220 22350 -40140 22360
rect -40220 22310 -40210 22350
rect -40710 22290 -40210 22310
rect -40150 22290 -40140 22350
rect -38690 22310 -38680 22370
rect -38620 22330 -38610 22370
rect -38500 22340 -38490 22400
rect -38430 22340 -38420 22400
rect -38500 22330 -38420 22340
rect -38130 22370 -38050 22380
rect -38130 22330 -38120 22370
rect -38620 22310 -38120 22330
rect -38060 22310 -38050 22370
rect -38690 22300 -38050 22310
rect -40780 22280 -40140 22290
rect -38320 22070 -38240 22080
rect -40480 22050 -40400 22060
rect -40780 22020 -40700 22030
rect -40780 21960 -40770 22020
rect -40710 21980 -40700 22020
rect -40480 21990 -40470 22050
rect -40410 21990 -40400 22050
rect -38690 22040 -38610 22050
rect -40480 21980 -40400 21990
rect -40220 22020 -40140 22030
rect -40220 21980 -40210 22020
rect -40710 21960 -40210 21980
rect -40150 21960 -40140 22020
rect -38690 21980 -38680 22040
rect -38620 22000 -38610 22040
rect -38320 22010 -38310 22070
rect -38250 22010 -38240 22070
rect -38320 22000 -38240 22010
rect -38130 22040 -38050 22050
rect -38130 22000 -38120 22040
rect -38620 21980 -38120 22000
rect -38060 21980 -38050 22040
rect -38690 21970 -38050 21980
rect -40780 21950 -40140 21960
rect -35940 21460 -35910 23210
rect -36130 21450 -35910 21460
rect -36130 21390 -36120 21450
rect -36060 21430 -35910 21450
rect -36060 21390 -36050 21430
rect -36130 21380 -36050 21390
rect -38500 20160 -38420 20170
rect -40590 20140 -40510 20150
rect -40780 20110 -40700 20120
rect -40780 20050 -40770 20110
rect -40710 20070 -40700 20110
rect -40590 20080 -40580 20140
rect -40520 20080 -40510 20140
rect -38690 20130 -38610 20140
rect -40590 20070 -40510 20080
rect -40220 20110 -40140 20120
rect -40220 20070 -40210 20110
rect -40710 20050 -40210 20070
rect -40150 20050 -40140 20110
rect -38690 20070 -38680 20130
rect -38620 20090 -38610 20130
rect -38500 20100 -38490 20160
rect -38430 20100 -38420 20160
rect -38500 20090 -38420 20100
rect -38130 20130 -38050 20140
rect -38130 20090 -38120 20130
rect -38620 20070 -38120 20090
rect -38060 20070 -38050 20130
rect -38690 20060 -38050 20070
rect -40780 20040 -40140 20050
rect -38320 19830 -38240 19840
rect -40480 19800 -40400 19810
rect -40780 19770 -40700 19780
rect -40780 19710 -40770 19770
rect -40710 19730 -40700 19770
rect -40480 19740 -40470 19800
rect -40410 19740 -40400 19800
rect -38690 19800 -38610 19810
rect -40480 19730 -40400 19740
rect -40220 19770 -40140 19780
rect -40220 19730 -40210 19770
rect -40710 19710 -40210 19730
rect -40150 19710 -40140 19770
rect -38690 19740 -38680 19800
rect -38620 19760 -38610 19800
rect -38320 19770 -38310 19830
rect -38250 19770 -38240 19830
rect -38320 19760 -38240 19770
rect -38130 19800 -38050 19810
rect -38130 19760 -38120 19800
rect -38620 19740 -38120 19760
rect -38060 19740 -38050 19800
rect -38690 19730 -38050 19740
rect -40780 19700 -40140 19710
rect -36120 19680 -36040 19690
rect -36120 19620 -36110 19680
rect -36050 19640 -36040 19680
rect -35940 19640 -35910 21430
rect -36050 19620 -35910 19640
rect -36120 19610 -35910 19620
rect -35940 19250 -35910 19610
rect -36120 19240 -35910 19250
rect -36120 19180 -36110 19240
rect -36050 19220 -35910 19240
rect -36050 19180 -36040 19220
rect -36120 19170 -36040 19180
rect -37700 18390 -37620 18400
rect -37700 18330 -37690 18390
rect -37630 18330 -37620 18390
rect -37700 18320 -37620 18330
rect -37700 18190 -37670 18320
rect -37700 18180 -37620 18190
rect -37700 18120 -37690 18180
rect -37630 18120 -37620 18180
rect -37700 18110 -37620 18120
rect -40590 17980 -40510 17990
rect -40590 17920 -40580 17980
rect -40520 17920 -40510 17980
rect -40590 17910 -40510 17920
rect -40590 17750 -40560 17910
rect -40590 17740 -40510 17750
rect -40590 17680 -40580 17740
rect -40520 17680 -40510 17740
rect -40590 17670 -40510 17680
rect -35940 17510 -35910 19220
rect -36120 17500 -35910 17510
rect -36120 17440 -36110 17500
rect -36050 17480 -35910 17500
rect -36050 17440 -36040 17480
rect -36120 17430 -36040 17440
rect -40590 17240 -40510 17250
rect -40590 17180 -40580 17240
rect -40520 17180 -40510 17240
rect -40590 17170 -40510 17180
rect -38580 17210 -38500 17220
rect -40590 17080 -40560 17170
rect -38580 17150 -38570 17210
rect -38510 17170 -38500 17210
rect -38210 17210 -38130 17220
rect -38210 17170 -38200 17210
rect -38510 17150 -38200 17170
rect -38140 17150 -38130 17210
rect -38580 17140 -38130 17150
rect -35940 17080 -35910 17480
rect -40590 17070 -40510 17080
rect -40590 17010 -40580 17070
rect -40520 17010 -40510 17070
rect -40590 17000 -40510 17010
rect -36120 17070 -35910 17080
rect -36120 17010 -36110 17070
rect -36050 17050 -35910 17070
rect -36050 17010 -36040 17050
rect -36120 17000 -36040 17010
rect -39990 15220 -39910 15230
rect -39990 15160 -39980 15220
rect -39920 15190 -39910 15220
rect -39920 15180 -39490 15190
rect -39920 15160 -39560 15180
rect -39990 15150 -39910 15160
rect -39570 15120 -39560 15160
rect -39500 15120 -39490 15180
rect -39570 15110 -39490 15120
rect -36190 14900 -36110 14910
rect -36190 14840 -36180 14900
rect -36120 14840 -36110 14900
rect -36190 14830 -36110 14840
rect -35220 10700 -35110 10720
rect -35220 10630 -35200 10700
rect -35130 10630 -35110 10700
rect -35220 10610 -35110 10630
rect -33810 10510 -33780 23260
rect -33600 18840 -33570 23320
rect -27200 23340 -27120 23350
rect -27200 23280 -27190 23340
rect -27130 23280 -27120 23340
rect -27200 23270 -27120 23280
rect -29440 21570 -29360 21580
rect -29440 21510 -29430 21570
rect -29370 21510 -29360 21570
rect -29440 21500 -29360 21510
rect -33600 18810 -32200 18840
rect -32230 18140 -32200 18810
rect -29440 18200 -29410 21500
rect -29380 20700 -27380 20710
rect -29380 20640 -29370 20700
rect -29310 20680 -27450 20700
rect -29310 20640 -29300 20680
rect -29380 20630 -29300 20640
rect -27460 20640 -27450 20680
rect -27390 20640 -27380 20700
rect -27460 20630 -27380 20640
rect -28390 18570 -28310 18580
rect -28390 18530 -28380 18570
rect -28450 18510 -28380 18530
rect -28320 18510 -28310 18570
rect -28450 18500 -28310 18510
rect -28450 18240 -28420 18500
rect -28390 18450 -28310 18460
rect -28390 18390 -28380 18450
rect -28320 18390 -28310 18450
rect -28390 18380 -28310 18390
rect -28340 18240 -28310 18380
rect -32120 18170 -29410 18200
rect -28500 18230 -28420 18240
rect -28500 18170 -28490 18230
rect -28430 18170 -28420 18230
rect -32230 18130 -32150 18140
rect -32230 18070 -32220 18130
rect -32160 18070 -32150 18130
rect -32230 18060 -32150 18070
rect -32120 17960 -32090 18170
rect -28500 18160 -28420 18170
rect -28390 18230 -28310 18240
rect -28390 18170 -28380 18230
rect -28320 18170 -28310 18230
rect -28390 18160 -28310 18170
rect -32060 18130 -31980 18140
rect -32060 18070 -32050 18130
rect -31990 18090 -31980 18130
rect -31990 18070 -24510 18090
rect -32060 18060 -24510 18070
rect -32170 17950 -32090 17960
rect -32170 17890 -32160 17950
rect -32100 17890 -32090 17950
rect -32170 17880 -32090 17890
rect -28630 17900 -28550 17910
rect -28630 17840 -28620 17900
rect -28560 17860 -28550 17900
rect -28210 17900 -28130 17910
rect -28210 17860 -28200 17900
rect -28560 17840 -28200 17860
rect -28140 17840 -28130 17900
rect -28630 17830 -28130 17840
rect -24540 17720 -24510 18060
rect -24540 17690 -22450 17720
rect -28390 17510 -28310 17520
rect -28390 17470 -28380 17510
rect -28580 17450 -28380 17470
rect -28320 17450 -28310 17510
rect -28580 17440 -28310 17450
rect -28580 17410 -28550 17440
rect -28630 17400 -28550 17410
rect -28630 17340 -28620 17400
rect -28560 17340 -28550 17400
rect -28630 17330 -28550 17340
rect -28450 17400 -28370 17410
rect -28450 17340 -28440 17400
rect -28380 17360 -28370 17400
rect -28210 17400 -28130 17410
rect -28210 17360 -28200 17400
rect -28380 17340 -28200 17360
rect -28140 17340 -28130 17400
rect -28450 17330 -28130 17340
rect -23990 17380 -23960 17690
rect -23270 17380 -23240 17690
rect -23990 17370 -23910 17380
rect -23990 17310 -23980 17370
rect -23920 17310 -23910 17370
rect -23990 17300 -23910 17310
rect -23270 17370 -23190 17380
rect -23270 17310 -23260 17370
rect -23200 17310 -23190 17370
rect -23270 17300 -23190 17310
rect -22480 16050 -22450 17690
rect -22480 16040 -22290 16050
rect -22480 16020 -22360 16040
rect -22370 15980 -22360 16020
rect -22300 15980 -22290 16040
rect -22370 15970 -22290 15980
rect -21950 15860 -21870 15870
rect -21950 15800 -21940 15860
rect -21880 15820 -21870 15860
rect -21770 15860 -21690 15870
rect -21770 15820 -21760 15860
rect -21880 15800 -21760 15820
rect -21700 15800 -21690 15860
rect -21950 15790 -21690 15800
rect -22620 15580 -22540 15590
rect -22970 15530 -22890 15540
rect -22970 15470 -22960 15530
rect -22900 15470 -22890 15530
rect -22620 15520 -22610 15580
rect -22550 15520 -22540 15580
rect -22620 15510 -22540 15520
rect -22970 15460 -22890 15470
rect -24530 15430 -24450 15440
rect -24530 15370 -24520 15430
rect -24460 15420 -24450 15430
rect -24460 15410 -24270 15420
rect -24460 15390 -24340 15410
rect -24460 15370 -24450 15390
rect -24530 15360 -24450 15370
rect -24350 15350 -24340 15390
rect -24280 15350 -24270 15410
rect -24350 15340 -24270 15350
rect -23810 15260 -23730 15270
rect -23810 15230 -23800 15260
rect -24480 15200 -23800 15230
rect -23740 15230 -23730 15260
rect -23270 15260 -23190 15270
rect -23270 15230 -23260 15260
rect -23740 15200 -23260 15230
rect -23200 15200 -23190 15260
rect -28620 14240 -28540 14250
rect -28620 14180 -28610 14240
rect -28550 14200 -28540 14240
rect -28220 14240 -28140 14250
rect -28220 14200 -28210 14240
rect -28550 14180 -28210 14200
rect -28150 14180 -28140 14240
rect -28620 14170 -28140 14180
rect -28630 13740 -28550 13750
rect -28630 13680 -28620 13740
rect -28560 13700 -28550 13740
rect -28210 13740 -28130 13750
rect -28210 13700 -28200 13740
rect -28560 13680 -28200 13700
rect -28140 13680 -28130 13740
rect -28630 13670 -28130 13680
rect -28630 13340 -28130 13350
rect -28630 13280 -28620 13340
rect -28560 13320 -28200 13340
rect -28560 13280 -28550 13320
rect -28630 13270 -28550 13280
rect -28210 13280 -28200 13320
rect -28140 13280 -28130 13340
rect -28210 13270 -28130 13280
rect -28630 13220 -28550 13230
rect -28630 13160 -28620 13220
rect -28560 13180 -28550 13220
rect -28210 13220 -28130 13230
rect -28210 13180 -28200 13220
rect -28560 13160 -28200 13180
rect -28140 13160 -28130 13220
rect -28630 13150 -28130 13160
rect -24480 12730 -24450 15200
rect -23810 15190 -23730 15200
rect -23270 15190 -23190 15200
rect -22970 15210 -22940 15460
rect -22570 15230 -22540 15510
rect -21770 15230 -21740 15790
rect -22970 15200 -22890 15210
rect -22570 15200 -21740 15230
rect -22970 15140 -22960 15200
rect -22900 15140 -22890 15200
rect -22970 15130 -22890 15140
rect -28630 12720 -28550 12730
rect -28630 12660 -28620 12720
rect -28560 12680 -28550 12720
rect -28450 12720 -28370 12730
rect -28450 12680 -28440 12720
rect -28560 12660 -28440 12680
rect -28380 12660 -28370 12720
rect -28630 12650 -28370 12660
rect -24600 12720 -24450 12730
rect -24600 12660 -24590 12720
rect -24530 12700 -24450 12720
rect -24530 12660 -24520 12700
rect -24600 12650 -24520 12660
rect -35220 10480 -33780 10510
rect -35220 8720 -35180 10480
rect -28620 9560 -28540 9570
rect -28620 9500 -28610 9560
rect -28550 9520 -28540 9560
rect -28220 9560 -28140 9570
rect -28220 9520 -28210 9560
rect -28550 9500 -28210 9520
rect -28150 9500 -28140 9560
rect -28620 9490 -28140 9500
rect -28630 9060 -28130 9070
rect -28630 9000 -28620 9060
rect -28560 9040 -28200 9060
rect -28560 9000 -28550 9040
rect -28630 8990 -28550 9000
rect -28210 9000 -28200 9040
rect -28140 9000 -28130 9060
rect -28210 8990 -28130 9000
rect -35260 8710 -35180 8720
rect -35260 8650 -35250 8710
rect -35190 8650 -35180 8710
rect -35260 8640 -35180 8650
rect -28620 8600 -28140 8610
rect -28620 8540 -28610 8600
rect -28550 8580 -28210 8600
rect -28550 8540 -28540 8580
rect -28620 8530 -28540 8540
rect -28220 8540 -28210 8580
rect -28150 8540 -28140 8600
rect -28220 8530 -28140 8540
rect -28390 8150 -28310 8160
rect -28390 8110 -28380 8150
rect -28580 8090 -28380 8110
rect -28320 8090 -28310 8150
rect -28580 8080 -28310 8090
rect -28580 8050 -28550 8080
rect -28630 8040 -28550 8050
rect -28630 7980 -28620 8040
rect -28560 7980 -28550 8040
rect -28630 7970 -28550 7980
rect -28450 8040 -28370 8050
rect -28450 7980 -28440 8040
rect -28380 8000 -28370 8040
rect -28210 8040 -28130 8050
rect -28210 8000 -28200 8040
rect -28380 7980 -28200 8000
rect -28140 7980 -28130 8040
rect -28450 7970 -28130 7980
rect -28620 4860 -28140 4870
rect -28620 4800 -28610 4860
rect -28550 4840 -28210 4860
rect -28550 4800 -28540 4840
rect -28620 4790 -28540 4800
rect -28220 4800 -28210 4840
rect -28150 4800 -28140 4860
rect -28220 4790 -28140 4800
rect -28560 4360 -28480 4370
rect -28560 4300 -28550 4360
rect -28490 4300 -28480 4360
rect -28560 4290 -28480 4300
rect -28280 4360 -28200 4370
rect -28280 4300 -28270 4360
rect -28210 4300 -28200 4360
rect -28280 4290 -28200 4300
rect -28280 4170 -28250 4290
rect -28620 4140 -28250 4170
rect -35150 4030 -35040 4050
rect -35150 3960 -35130 4030
rect -35060 3960 -35040 4030
rect -35150 3940 -35040 3960
rect -28620 3850 -28590 4140
rect -28560 4100 -28480 4110
rect -28560 4040 -28550 4100
rect -28490 4040 -28480 4100
rect -28560 4030 -28480 4040
rect -28510 4000 -28480 4030
rect -28510 3970 -28250 4000
rect -28280 3850 -28250 3970
rect -28620 3840 -28480 3850
rect -28620 3820 -28550 3840
rect -28560 3780 -28550 3820
rect -28490 3780 -28480 3840
rect -28560 3770 -28480 3780
rect -28280 3840 -28200 3850
rect -28280 3780 -28270 3840
rect -28210 3780 -28200 3840
rect -28280 3770 -28200 3780
rect -21700 3510 -21620 3520
rect -28390 3450 -28310 3460
rect -28390 3390 -28380 3450
rect -28320 3390 -28310 3450
rect -21700 3450 -21690 3510
rect -21630 3450 -21620 3510
rect -21700 3440 -21620 3450
rect -28390 3380 -28310 3390
rect -28630 3340 -28550 3350
rect -28630 3280 -28620 3340
rect -28560 3300 -28550 3340
rect -28450 3340 -28370 3350
rect -28450 3300 -28440 3340
rect -28560 3280 -28440 3300
rect -28380 3280 -28370 3340
rect -28630 3270 -28370 3280
rect -28340 3300 -28310 3380
rect -21650 3350 -21620 3440
rect -28210 3340 -28130 3350
rect -28210 3300 -28200 3340
rect -28340 3280 -28200 3300
rect -28140 3280 -28130 3340
rect -28340 3270 -28130 3280
rect -21700 3340 -21620 3350
rect -21700 3280 -21690 3340
rect -21630 3280 -21620 3340
rect -21700 3270 -21620 3280
rect -28620 160 -28140 170
rect -28620 100 -28610 160
rect -28550 140 -28210 160
rect -28550 100 -28540 140
rect -28620 90 -28540 100
rect -28220 100 -28210 140
rect -28150 100 -28140 160
rect -28220 90 -28140 100
rect -28620 -400 -28540 -390
rect -28620 -460 -28610 -400
rect -28550 -440 -28540 -400
rect -28220 -400 -28140 -390
rect -28220 -440 -28210 -400
rect -28550 -460 -28210 -440
rect -28150 -460 -28140 -400
rect -28620 -470 -28140 -460
rect -28590 -600 -28480 -580
rect -28590 -670 -28570 -600
rect -28500 -670 -28480 -600
rect -28590 -690 -28480 -670
rect -28390 -600 -28280 -580
rect -28390 -670 -28370 -600
rect -28300 -670 -28280 -600
rect -28390 -690 -28280 -670
rect -15000 -730 -14890 -710
rect -15000 -800 -14980 -730
rect -14910 -800 -14890 -730
rect -15000 -820 -14890 -800
<< via2 >>
rect -26660 24680 -26590 24750
rect -21330 24780 -21260 24850
rect -21000 24750 -20930 24820
rect -35200 10630 -35130 10700
rect -35130 3960 -35060 4030
rect -28570 -670 -28500 -600
rect -28370 -670 -28300 -600
rect -14980 -800 -14910 -730
<< metal3 >>
rect -21350 24850 -21240 24870
rect -21350 24780 -21330 24850
rect -21260 24780 -21240 24850
rect -26680 24750 -26570 24770
rect -21350 24760 -21240 24780
rect -21020 24820 -20910 24840
rect -26680 24680 -26660 24750
rect -26590 24680 -26570 24750
rect -21020 24750 -21000 24820
rect -20930 24750 -20910 24820
rect -21020 24730 -20910 24750
rect -26680 24660 -26570 24680
rect -35220 10700 -35110 10720
rect -35220 10630 -35200 10700
rect -35130 10630 -35110 10700
rect -35220 10610 -35110 10630
rect -35150 4030 -35040 4050
rect -35150 3960 -35130 4030
rect -35060 3960 -35040 4030
rect -35150 3940 -35040 3960
rect -28590 -600 -28480 -580
rect -28590 -670 -28570 -600
rect -28500 -670 -28480 -600
rect -28590 -690 -28480 -670
rect -28390 -600 -28280 -580
rect -28390 -670 -28370 -600
rect -28300 -670 -28280 -600
rect -28390 -690 -28280 -670
rect -15000 -730 -14890 -710
rect -15000 -800 -14980 -730
rect -14910 -800 -14890 -730
rect -15000 -820 -14890 -800
<< via3 >>
rect -21330 24780 -21260 24850
rect -26660 24680 -26590 24750
rect -21000 24750 -20930 24820
rect -35200 10630 -35130 10700
rect -35130 3960 -35060 4030
rect -28570 -670 -28500 -600
rect -28370 -670 -28300 -600
rect -14980 -800 -14910 -730
<< metal4 >>
rect -26600 27250 -26540 27650
rect -20930 27500 -20790 27650
rect -26600 24770 -26540 25330
rect -26680 24750 -26540 24770
rect -21350 24850 -21240 24870
rect -21350 24780 -21330 24850
rect -21260 24780 -21240 24850
rect -21010 24840 -20910 25280
rect -21350 24760 -21240 24780
rect -26680 24680 -26660 24750
rect -26590 24680 -26540 24750
rect -26680 24660 -26540 24680
rect -26600 18180 -26540 24660
rect -21300 24670 -21240 24760
rect -21020 24820 -20910 24840
rect -21020 24750 -21000 24820
rect -20930 24750 -20910 24820
rect -21020 24730 -20910 24750
rect -20850 24670 -20790 27500
rect -21300 24610 -20790 24670
rect -26600 18120 -24420 18180
rect -24480 17810 -24420 18120
rect -24480 17750 -22360 17810
rect -22420 16220 -22360 17750
rect -22420 16160 -20680 16220
rect -35220 10700 -35110 10720
rect -35220 10670 -35200 10700
rect -35740 10630 -35200 10670
rect -35130 10630 -35110 10700
rect -35740 10610 -35110 10630
rect -35740 10470 -35680 10610
rect -20740 10470 -20680 16160
rect -41600 4740 -41540 5150
rect -35390 4800 -35330 5100
rect -21360 4740 -21300 5150
rect -15170 4790 -15070 5090
rect -35150 4030 -35040 4050
rect -35150 4000 -35130 4030
rect -35330 3960 -35130 4000
rect -35060 3960 -35040 4030
rect -35330 3940 -35040 3960
rect -21550 -380 -21360 -360
rect -22150 -420 -21360 -380
rect -41600 -970 -41540 -420
rect -22150 -440 -21490 -420
rect -35400 -500 -35310 -470
rect -35400 -560 -28710 -500
rect -35400 -910 -35320 -560
rect -28910 -620 -28710 -560
rect -28590 -600 -28480 -580
rect -28590 -670 -28570 -600
rect -28500 -670 -28480 -600
rect -28590 -690 -28480 -670
rect -28390 -600 -28280 -580
rect -28390 -670 -28370 -600
rect -28300 -670 -28280 -600
rect -28390 -690 -28280 -670
rect -22150 -680 -21950 -440
rect -21760 -660 -21520 -500
rect -22100 -720 -21950 -680
rect -21630 -670 -21520 -660
rect -15170 -670 -15070 -480
rect -21630 -710 -15070 -670
rect -21630 -730 -14890 -710
rect -15170 -800 -14980 -730
rect -14910 -800 -14890 -730
rect -15170 -820 -14890 -800
rect -15170 -920 -15070 -820
rect -35750 -6420 -35690 -5990
rect -35100 -6420 -34930 -5930
rect -22150 -6080 -21950 -5990
rect -22010 -6130 -21950 -6080
rect -21360 -6130 -21300 -5990
rect -22010 -6190 -21300 -6130
rect -35750 -6480 -34930 -6420
use bias_generator  bias_generator_0
timestamp 1730563144
transform 1 0 -44836 0 1 8370
box 3156 2360 10700 6640
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_0
timestamp 1730563144
transform 1 0 -31884 0 1 -3330
box -3186 -2740 3186 2740
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_1
timestamp 1730563144
transform 1 0 -38504 0 1 -3630
box -3186 -2740 3186 2740
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_2
timestamp 1730563144
transform 1 0 -38504 0 1 2090
box -3186 -2740 3186 2740
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_3
timestamp 1730563144
transform 1 0 -18254 0 1 2090
box -3186 -2740 3186 2740
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_4
timestamp 1730563144
transform 1 0 -24900 0 1 -3334
box -3186 -2740 3186 2740
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_5
timestamp 1730563144
transform 1 0 -18254 0 1 -3630
box -3186 -2740 3186 2740
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  sky130_fd_pr__cap_mim_m3_1_5HBWYY_6
timestamp 1730563144
transform 1 0 -18254 0 1 7810
box -3186 -2740 3186 2740
use sky130_fd_pr__nfet_01v8_lvt_C84B7J  sky130_fd_pr__nfet_01v8_lvt_C84B7J_0
timestamp 1730563144
transform 1 0 -27954 0 1 21239
box -296 -379 296 379
use sky130_fd_pr__nfet_01v8_lvt_FWQUH5  sky130_fd_pr__nfet_01v8_lvt_FWQUH5_0
timestamp 1730563144
transform 1 0 -36534 0 1 18340
box -596 -1010 596 1010
use sky130_fd_pr__nfet_01v8_lvt_N28DAC  sky130_fd_pr__nfet_01v8_lvt_N28DAC_0
timestamp 1730563144
transform 1 0 -32884 0 1 9210
box -596 -510 596 510
use sky130_fd_pr__nfet_01v8_lvt_Q53FMB  sky130_fd_pr__nfet_01v8_lvt_Q53FMB_0
timestamp 1730563144
transform 1 0 -31109 0 1 24300
box -231 -460 231 460
use sky130_fd_pr__nfet_01v8_lvt_QW8YAA  sky130_fd_pr__nfet_01v8_lvt_QW8YAA_0
timestamp 1730563144
transform 1 0 -30335 0 1 15790
box -1825 -2210 1825 2210
use sky130_fd_pr__nfet_01v8_lvt_QW8YAA  sky130_fd_pr__nfet_01v8_lvt_QW8YAA_1
timestamp 1730563144
transform 1 0 -30335 0 1 11110
box -1825 -2210 1825 2210
use sky130_fd_pr__nfet_01v8_lvt_QW8YAA  sky130_fd_pr__nfet_01v8_lvt_QW8YAA_2
timestamp 1730563144
transform 1 0 -22625 0 1 12920
box -1825 -2210 1825 2210
use sky130_fd_pr__nfet_01v8_lvt_SHAVFW  sky130_fd_pr__nfet_01v8_lvt_SHAVFW_0
timestamp 1730563144
transform 1 0 -28335 0 1 23949
box -1255 -819 1255 819
use sky130_fd_pr__nfet_01v8_lvt_W9NHZX  sky130_fd_pr__nfet_01v8_lvt_W9NHZX_0
timestamp 1730563144
transform 1 0 -37459 0 1 17790
box -231 -460 231 460
use sky130_fd_pr__nfet_01v8_lvt_W9NHZX  sky130_fd_pr__nfet_01v8_lvt_W9NHZX_1
timestamp 1730563144
transform 1 0 -37459 0 1 15620
box -231 -460 231 460
use sky130_fd_pr__nfet_01v8_lvt_WA2NKZ  sky130_fd_pr__nfet_01v8_lvt_WA2NKZ_0
timestamp 1730563144
transform 1 0 -34414 0 1 19201
box -596 -4191 596 4191
use sky130_fd_pr__pfet_01v8_JHT74A  sky130_fd_pr__pfet_01v8_JHT74A_0
timestamp 1730563144
transform 1 0 -27885 0 1 19459
box -365 -1219 365 1219
use sky130_fd_pr__pfet_01v8_lvt_545GKL  sky130_fd_pr__pfet_01v8_lvt_545GKL_0
timestamp 1730563144
transform 1 0 -31845 0 1 6419
box -3335 -2219 3335 2219
use sky130_fd_pr__pfet_01v8_lvt_545GKL  sky130_fd_pr__pfet_01v8_lvt_545GKL_1
timestamp 1730563144
transform 1 0 -24915 0 1 6419
box -3335 -2219 3335 2219
use sky130_fd_pr__pfet_01v8_lvt_545GKL  sky130_fd_pr__pfet_01v8_lvt_545GKL_2
timestamp 1730563144
transform 1 0 -31845 0 1 1719
box -3335 -2219 3335 2219
use sky130_fd_pr__pfet_01v8_lvt_MF6SRL  sky130_fd_pr__pfet_01v8_lvt_MF6SRL_0
timestamp 1730563144
transform 1 0 -38009 0 1 22343
box -231 -4573 231 4573
use sky130_fd_pr__pfet_01v8_lvt_MXC9RL  sky130_fd_pr__pfet_01v8_lvt_MXC9RL_0
timestamp 1730563144
transform 1 0 -33829 0 1 25927
box -231 -2337 231 2337
use sky130_fd_pr__pfet_01v8_M5XJZ4  sky130_fd_pr__pfet_01v8_M5XJZ4_0
timestamp 1730563144
transform 1 0 -41146 0 1 28359
box -554 -1219 554 1219
use sky130_fd_pr__pfet_01v8_M7ZEKL  sky130_fd_pr__pfet_01v8_M7ZEKL_0
timestamp 1730563144
transform 1 0 -22779 0 1 16449
box -231 -1219 231 1219
use sky130_fd_pr__pfet_01v8_MD8735  sky130_fd_pr__pfet_01v8_MD8735_0
timestamp 1730563144
transform 1 0 -34876 0 1 25927
box -554 -2337 554 2337
use sky130_fd_pr__pfet_01v8_MV5GT4  sky130_fd_pr__pfet_01v8_MV5GT4_0
timestamp 1730563144
transform 1 0 -39056 0 1 22343
box -554 -4573 554 4573
use sky130_fd_pr__cap_mim_m3_1_A4BC7Z  XC1
timestamp 1730563144
transform 1 0 -23794 0 1 26290
box -2886 -1040 2886 1040
use sky130_fd_pr__cap_mim_m3_1_A4BC7Z  XC2
timestamp 1730563144
transform 1 0 -23794 0 1 28610
box -2886 -1040 2886 1040
use sky130_fd_pr__cap_mim_m3_1_5HBWYY  XC3
timestamp 1730563144
transform 1 0 -38494 0 1 7810
box -3186 -2740 3186 2740
use sky130_fd_pr__pfet_01v8_lvt_QQJVLQ  XM2
timestamp 1730563144
transform 1 0 -28339 0 1 27217
box -871 -2337 871 2337
use sky130_fd_pr__nfet_01v8_lvt_Q53FMB  XM4
timestamp 1730563144
transform 1 0 -30379 0 1 24310
box -231 -460 231 460
use sky130_fd_pr__nfet_01v8_lvt_Q53FMB  XM5
timestamp 1730563144
transform 1 0 -31829 0 1 24300
box -231 -460 231 460
use sky130_fd_pr__pfet_01v8_lvt_PD3USF  XM6
timestamp 1730563144
transform 1 0 -30379 0 1 28339
box -231 -1219 231 1219
use sky130_fd_pr__pfet_01v8_lvt_SLP2FE  XM7
timestamp 1730563144
transform 1 0 -31099 0 1 28339
box -231 -1219 231 1219
use sky130_fd_pr__pfet_01v8_lvt_SLP2FE  XM8
timestamp 1730563144
transform 1 0 -31819 0 1 28339
box -231 -1219 231 1219
use sky130_fd_pr__nfet_01v8_lvt_C84B7J  XM10
timestamp 1730563144
transform 1 0 -28804 0 1 21239
box -296 -379 296 379
use sky130_fd_pr__pfet_01v8_JHT74A  XM11
timestamp 1730563144
transform 1 0 -28875 0 1 19459
box -365 -1219 365 1219
use sky130_fd_pr__nfet_01v8_lvt_QW8YAA  XM13
timestamp 1730563144
transform 1 0 -26425 0 1 11110
box -1825 -2210 1825 2210
use sky130_fd_pr__nfet_01v8_lvt_QW8YAA  XM14
timestamp 1730563144
transform 1 0 -26425 0 1 15790
box -1825 -2210 1825 2210
use sky130_fd_pr__pfet_01v8_lvt_545GKL  XM16
timestamp 1730563144
transform 1 0 -24915 0 1 1719
box -3335 -2219 3335 2219
use sky130_fd_pr__pfet_01v8_M7ZEKL  XM17
timestamp 1730563144
transform 1 0 -24219 0 1 16449
box -231 -1219 231 1219
use sky130_fd_pr__pfet_01v8_M7ZEKL  XM18
timestamp 1730563144
transform 1 0 -23499 0 1 16449
box -231 -1219 231 1219
use sky130_fd_pr__nfet_01v8_lvt_N28DAC  XM21
timestamp 1730563144
transform 1 0 -34164 0 1 9210
box -596 -510 596 510
use sky130_fd_pr__nfet_01v8_lvt_WA2NKZ  XM24
timestamp 1730563144
transform 1 0 -32884 0 1 14441
box -596 -4191 596 4191
use sky130_fd_pr__pfet_01v8_M5XJZ4  XM25
timestamp 1730563144
transform 1 0 -39056 0 1 16289
box -554 -1219 554 1219
use sky130_fd_pr__pfet_01v8_M5XJZ4  XM26
timestamp 1730563144
transform 1 0 -41146 0 1 16259
box -554 -1219 554 1219
use sky130_fd_pr__pfet_01v8_lvt_M7ZRRL  XM27
timestamp 1730563144
transform 1 0 -38009 0 1 16289
box -231 -1219 231 1219
use sky130_fd_pr__pfet_01v8_lvt_M7ZRRL  XM28
timestamp 1730563144
transform 1 0 -40099 0 1 16259
box -231 -1219 231 1219
use sky130_fd_pr__nfet_01v8_lvt_FWQUH5  XM31
timestamp 1730563144
transform 1 0 -36533 0 1 16171
box -596 -1010 596 1010
use sky130_fd_pr__nfet_01v8_lvt_PP2UM9  XM34
timestamp 1730563144
transform 1 0 -36534 0 1 21419
box -596 -1919 596 1919
use sky130_fd_pr__pfet_01v8_lvt_M7ZRRL  XM35
timestamp 1730563144
transform 1 0 -40099 0 1 28359
box -231 -1219 231 1219
use sky130_fd_pr__pfet_01v8_MD8735  XM36
timestamp 1730563144
transform 1 0 -36966 0 1 25927
box -554 -2337 554 2337
use sky130_fd_pr__pfet_01v8_lvt_MXC9RL  XM37
timestamp 1730563144
transform 1 0 -35919 0 1 25927
box -231 -2337 231 2337
use sky130_fd_pr__pfet_01v8_MV5GT4  XM40
timestamp 1730563144
transform 1 0 -41146 0 1 22313
box -554 -4573 554 4573
use sky130_fd_pr__pfet_01v8_lvt_MF6SRL  XM41
timestamp 1730563144
transform 1 0 -40099 0 1 22313
box -231 -4573 231 4573
use sky130_fd_pr__pfet_01v8_F4HV3A  XM44
timestamp 1730563144
transform 1 0 -22059 0 1 15699
box -231 -469 231 469
<< end >>
