magic
tech sky130A
magscale 1 2
timestamp 1729530615
<< error_p >>
rect -1055 681 -993 687
rect -927 681 -865 687
rect -799 681 -737 687
rect -671 681 -609 687
rect -543 681 -481 687
rect -415 681 -353 687
rect -287 681 -225 687
rect -159 681 -97 687
rect -31 681 31 687
rect 97 681 159 687
rect 225 681 287 687
rect 353 681 415 687
rect 481 681 543 687
rect 609 681 671 687
rect 737 681 799 687
rect 865 681 927 687
rect 993 681 1055 687
rect -1055 647 -1043 681
rect -927 647 -915 681
rect -799 647 -787 681
rect -671 647 -659 681
rect -543 647 -531 681
rect -415 647 -403 681
rect -287 647 -275 681
rect -159 647 -147 681
rect -31 647 -19 681
rect 97 647 109 681
rect 225 647 237 681
rect 353 647 365 681
rect 481 647 493 681
rect 609 647 621 681
rect 737 647 749 681
rect 865 647 877 681
rect 993 647 1005 681
rect -1055 641 -993 647
rect -927 641 -865 647
rect -799 641 -737 647
rect -671 641 -609 647
rect -543 641 -481 647
rect -415 641 -353 647
rect -287 641 -225 647
rect -159 641 -97 647
rect -31 641 31 647
rect 97 641 159 647
rect 225 641 287 647
rect 353 641 415 647
rect 481 641 543 647
rect 609 641 671 647
rect 737 641 799 647
rect 865 641 927 647
rect 993 641 1055 647
rect -1055 71 -993 77
rect -927 71 -865 77
rect -799 71 -737 77
rect -671 71 -609 77
rect -543 71 -481 77
rect -415 71 -353 77
rect -287 71 -225 77
rect -159 71 -97 77
rect -31 71 31 77
rect 97 71 159 77
rect 225 71 287 77
rect 353 71 415 77
rect 481 71 543 77
rect 609 71 671 77
rect 737 71 799 77
rect 865 71 927 77
rect 993 71 1055 77
rect -1055 37 -1043 71
rect -927 37 -915 71
rect -799 37 -787 71
rect -671 37 -659 71
rect -543 37 -531 71
rect -415 37 -403 71
rect -287 37 -275 71
rect -159 37 -147 71
rect -31 37 -19 71
rect 97 37 109 71
rect 225 37 237 71
rect 353 37 365 71
rect 481 37 493 71
rect 609 37 621 71
rect 737 37 749 71
rect 865 37 877 71
rect 993 37 1005 71
rect -1055 31 -993 37
rect -927 31 -865 37
rect -799 31 -737 37
rect -671 31 -609 37
rect -543 31 -481 37
rect -415 31 -353 37
rect -287 31 -225 37
rect -159 31 -97 37
rect -31 31 31 37
rect 97 31 159 37
rect 225 31 287 37
rect 353 31 415 37
rect 481 31 543 37
rect 609 31 671 37
rect 737 31 799 37
rect 865 31 927 37
rect 993 31 1055 37
rect -1055 -37 -993 -31
rect -927 -37 -865 -31
rect -799 -37 -737 -31
rect -671 -37 -609 -31
rect -543 -37 -481 -31
rect -415 -37 -353 -31
rect -287 -37 -225 -31
rect -159 -37 -97 -31
rect -31 -37 31 -31
rect 97 -37 159 -31
rect 225 -37 287 -31
rect 353 -37 415 -31
rect 481 -37 543 -31
rect 609 -37 671 -31
rect 737 -37 799 -31
rect 865 -37 927 -31
rect 993 -37 1055 -31
rect -1055 -71 -1043 -37
rect -927 -71 -915 -37
rect -799 -71 -787 -37
rect -671 -71 -659 -37
rect -543 -71 -531 -37
rect -415 -71 -403 -37
rect -287 -71 -275 -37
rect -159 -71 -147 -37
rect -31 -71 -19 -37
rect 97 -71 109 -37
rect 225 -71 237 -37
rect 353 -71 365 -37
rect 481 -71 493 -37
rect 609 -71 621 -37
rect 737 -71 749 -37
rect 865 -71 877 -37
rect 993 -71 1005 -37
rect -1055 -77 -993 -71
rect -927 -77 -865 -71
rect -799 -77 -737 -71
rect -671 -77 -609 -71
rect -543 -77 -481 -71
rect -415 -77 -353 -71
rect -287 -77 -225 -71
rect -159 -77 -97 -71
rect -31 -77 31 -71
rect 97 -77 159 -71
rect 225 -77 287 -71
rect 353 -77 415 -71
rect 481 -77 543 -71
rect 609 -77 671 -71
rect 737 -77 799 -71
rect 865 -77 927 -71
rect 993 -77 1055 -71
rect -1055 -647 -993 -641
rect -927 -647 -865 -641
rect -799 -647 -737 -641
rect -671 -647 -609 -641
rect -543 -647 -481 -641
rect -415 -647 -353 -641
rect -287 -647 -225 -641
rect -159 -647 -97 -641
rect -31 -647 31 -641
rect 97 -647 159 -641
rect 225 -647 287 -641
rect 353 -647 415 -641
rect 481 -647 543 -641
rect 609 -647 671 -641
rect 737 -647 799 -641
rect 865 -647 927 -641
rect 993 -647 1055 -641
rect -1055 -681 -1043 -647
rect -927 -681 -915 -647
rect -799 -681 -787 -647
rect -671 -681 -659 -647
rect -543 -681 -531 -647
rect -415 -681 -403 -647
rect -287 -681 -275 -647
rect -159 -681 -147 -647
rect -31 -681 -19 -647
rect 97 -681 109 -647
rect 225 -681 237 -647
rect 353 -681 365 -647
rect 481 -681 493 -647
rect 609 -681 621 -647
rect 737 -681 749 -647
rect 865 -681 877 -647
rect 993 -681 1005 -647
rect -1055 -687 -993 -681
rect -927 -687 -865 -681
rect -799 -687 -737 -681
rect -671 -687 -609 -681
rect -543 -687 -481 -681
rect -415 -687 -353 -681
rect -287 -687 -225 -681
rect -159 -687 -97 -681
rect -31 -687 31 -681
rect 97 -687 159 -681
rect 225 -687 287 -681
rect 353 -687 415 -681
rect 481 -687 543 -681
rect 609 -687 671 -681
rect 737 -687 799 -681
rect 865 -687 927 -681
rect 993 -687 1055 -681
<< pwell >>
rect -1255 -819 1255 819
<< nmoslvt >>
rect -1059 109 -989 609
rect -931 109 -861 609
rect -803 109 -733 609
rect -675 109 -605 609
rect -547 109 -477 609
rect -419 109 -349 609
rect -291 109 -221 609
rect -163 109 -93 609
rect -35 109 35 609
rect 93 109 163 609
rect 221 109 291 609
rect 349 109 419 609
rect 477 109 547 609
rect 605 109 675 609
rect 733 109 803 609
rect 861 109 931 609
rect 989 109 1059 609
rect -1059 -609 -989 -109
rect -931 -609 -861 -109
rect -803 -609 -733 -109
rect -675 -609 -605 -109
rect -547 -609 -477 -109
rect -419 -609 -349 -109
rect -291 -609 -221 -109
rect -163 -609 -93 -109
rect -35 -609 35 -109
rect 93 -609 163 -109
rect 221 -609 291 -109
rect 349 -609 419 -109
rect 477 -609 547 -109
rect 605 -609 675 -109
rect 733 -609 803 -109
rect 861 -609 931 -109
rect 989 -609 1059 -109
<< ndiff >>
rect -1117 597 -1059 609
rect -1117 121 -1105 597
rect -1071 121 -1059 597
rect -1117 109 -1059 121
rect -989 597 -931 609
rect -989 121 -977 597
rect -943 121 -931 597
rect -989 109 -931 121
rect -861 597 -803 609
rect -861 121 -849 597
rect -815 121 -803 597
rect -861 109 -803 121
rect -733 597 -675 609
rect -733 121 -721 597
rect -687 121 -675 597
rect -733 109 -675 121
rect -605 597 -547 609
rect -605 121 -593 597
rect -559 121 -547 597
rect -605 109 -547 121
rect -477 597 -419 609
rect -477 121 -465 597
rect -431 121 -419 597
rect -477 109 -419 121
rect -349 597 -291 609
rect -349 121 -337 597
rect -303 121 -291 597
rect -349 109 -291 121
rect -221 597 -163 609
rect -221 121 -209 597
rect -175 121 -163 597
rect -221 109 -163 121
rect -93 597 -35 609
rect -93 121 -81 597
rect -47 121 -35 597
rect -93 109 -35 121
rect 35 597 93 609
rect 35 121 47 597
rect 81 121 93 597
rect 35 109 93 121
rect 163 597 221 609
rect 163 121 175 597
rect 209 121 221 597
rect 163 109 221 121
rect 291 597 349 609
rect 291 121 303 597
rect 337 121 349 597
rect 291 109 349 121
rect 419 597 477 609
rect 419 121 431 597
rect 465 121 477 597
rect 419 109 477 121
rect 547 597 605 609
rect 547 121 559 597
rect 593 121 605 597
rect 547 109 605 121
rect 675 597 733 609
rect 675 121 687 597
rect 721 121 733 597
rect 675 109 733 121
rect 803 597 861 609
rect 803 121 815 597
rect 849 121 861 597
rect 803 109 861 121
rect 931 597 989 609
rect 931 121 943 597
rect 977 121 989 597
rect 931 109 989 121
rect 1059 597 1117 609
rect 1059 121 1071 597
rect 1105 121 1117 597
rect 1059 109 1117 121
rect -1117 -121 -1059 -109
rect -1117 -597 -1105 -121
rect -1071 -597 -1059 -121
rect -1117 -609 -1059 -597
rect -989 -121 -931 -109
rect -989 -597 -977 -121
rect -943 -597 -931 -121
rect -989 -609 -931 -597
rect -861 -121 -803 -109
rect -861 -597 -849 -121
rect -815 -597 -803 -121
rect -861 -609 -803 -597
rect -733 -121 -675 -109
rect -733 -597 -721 -121
rect -687 -597 -675 -121
rect -733 -609 -675 -597
rect -605 -121 -547 -109
rect -605 -597 -593 -121
rect -559 -597 -547 -121
rect -605 -609 -547 -597
rect -477 -121 -419 -109
rect -477 -597 -465 -121
rect -431 -597 -419 -121
rect -477 -609 -419 -597
rect -349 -121 -291 -109
rect -349 -597 -337 -121
rect -303 -597 -291 -121
rect -349 -609 -291 -597
rect -221 -121 -163 -109
rect -221 -597 -209 -121
rect -175 -597 -163 -121
rect -221 -609 -163 -597
rect -93 -121 -35 -109
rect -93 -597 -81 -121
rect -47 -597 -35 -121
rect -93 -609 -35 -597
rect 35 -121 93 -109
rect 35 -597 47 -121
rect 81 -597 93 -121
rect 35 -609 93 -597
rect 163 -121 221 -109
rect 163 -597 175 -121
rect 209 -597 221 -121
rect 163 -609 221 -597
rect 291 -121 349 -109
rect 291 -597 303 -121
rect 337 -597 349 -121
rect 291 -609 349 -597
rect 419 -121 477 -109
rect 419 -597 431 -121
rect 465 -597 477 -121
rect 419 -609 477 -597
rect 547 -121 605 -109
rect 547 -597 559 -121
rect 593 -597 605 -121
rect 547 -609 605 -597
rect 675 -121 733 -109
rect 675 -597 687 -121
rect 721 -597 733 -121
rect 675 -609 733 -597
rect 803 -121 861 -109
rect 803 -597 815 -121
rect 849 -597 861 -121
rect 803 -609 861 -597
rect 931 -121 989 -109
rect 931 -597 943 -121
rect 977 -597 989 -121
rect 931 -609 989 -597
rect 1059 -121 1117 -109
rect 1059 -597 1071 -121
rect 1105 -597 1117 -121
rect 1059 -609 1117 -597
<< ndiffc >>
rect -1105 121 -1071 597
rect -977 121 -943 597
rect -849 121 -815 597
rect -721 121 -687 597
rect -593 121 -559 597
rect -465 121 -431 597
rect -337 121 -303 597
rect -209 121 -175 597
rect -81 121 -47 597
rect 47 121 81 597
rect 175 121 209 597
rect 303 121 337 597
rect 431 121 465 597
rect 559 121 593 597
rect 687 121 721 597
rect 815 121 849 597
rect 943 121 977 597
rect 1071 121 1105 597
rect -1105 -597 -1071 -121
rect -977 -597 -943 -121
rect -849 -597 -815 -121
rect -721 -597 -687 -121
rect -593 -597 -559 -121
rect -465 -597 -431 -121
rect -337 -597 -303 -121
rect -209 -597 -175 -121
rect -81 -597 -47 -121
rect 47 -597 81 -121
rect 175 -597 209 -121
rect 303 -597 337 -121
rect 431 -597 465 -121
rect 559 -597 593 -121
rect 687 -597 721 -121
rect 815 -597 849 -121
rect 943 -597 977 -121
rect 1071 -597 1105 -121
<< psubdiff >>
rect -1219 749 -1123 783
rect 1123 749 1219 783
rect -1219 687 -1185 749
rect 1185 687 1219 749
rect -1219 -749 -1185 -687
rect 1185 -749 1219 -687
rect -1219 -783 -1123 -749
rect 1123 -783 1219 -749
<< psubdiffcont >>
rect -1123 749 1123 783
rect -1219 -687 -1185 687
rect 1185 -687 1219 687
rect -1123 -783 1123 -749
<< poly >>
rect -1059 681 -989 697
rect -1059 647 -1043 681
rect -1005 647 -989 681
rect -1059 609 -989 647
rect -931 681 -861 697
rect -931 647 -915 681
rect -877 647 -861 681
rect -931 609 -861 647
rect -803 681 -733 697
rect -803 647 -787 681
rect -749 647 -733 681
rect -803 609 -733 647
rect -675 681 -605 697
rect -675 647 -659 681
rect -621 647 -605 681
rect -675 609 -605 647
rect -547 681 -477 697
rect -547 647 -531 681
rect -493 647 -477 681
rect -547 609 -477 647
rect -419 681 -349 697
rect -419 647 -403 681
rect -365 647 -349 681
rect -419 609 -349 647
rect -291 681 -221 697
rect -291 647 -275 681
rect -237 647 -221 681
rect -291 609 -221 647
rect -163 681 -93 697
rect -163 647 -147 681
rect -109 647 -93 681
rect -163 609 -93 647
rect -35 681 35 697
rect -35 647 -19 681
rect 19 647 35 681
rect -35 609 35 647
rect 93 681 163 697
rect 93 647 109 681
rect 147 647 163 681
rect 93 609 163 647
rect 221 681 291 697
rect 221 647 237 681
rect 275 647 291 681
rect 221 609 291 647
rect 349 681 419 697
rect 349 647 365 681
rect 403 647 419 681
rect 349 609 419 647
rect 477 681 547 697
rect 477 647 493 681
rect 531 647 547 681
rect 477 609 547 647
rect 605 681 675 697
rect 605 647 621 681
rect 659 647 675 681
rect 605 609 675 647
rect 733 681 803 697
rect 733 647 749 681
rect 787 647 803 681
rect 733 609 803 647
rect 861 681 931 697
rect 861 647 877 681
rect 915 647 931 681
rect 861 609 931 647
rect 989 681 1059 697
rect 989 647 1005 681
rect 1043 647 1059 681
rect 989 609 1059 647
rect -1059 71 -989 109
rect -1059 37 -1043 71
rect -1005 37 -989 71
rect -1059 21 -989 37
rect -931 71 -861 109
rect -931 37 -915 71
rect -877 37 -861 71
rect -931 21 -861 37
rect -803 71 -733 109
rect -803 37 -787 71
rect -749 37 -733 71
rect -803 21 -733 37
rect -675 71 -605 109
rect -675 37 -659 71
rect -621 37 -605 71
rect -675 21 -605 37
rect -547 71 -477 109
rect -547 37 -531 71
rect -493 37 -477 71
rect -547 21 -477 37
rect -419 71 -349 109
rect -419 37 -403 71
rect -365 37 -349 71
rect -419 21 -349 37
rect -291 71 -221 109
rect -291 37 -275 71
rect -237 37 -221 71
rect -291 21 -221 37
rect -163 71 -93 109
rect -163 37 -147 71
rect -109 37 -93 71
rect -163 21 -93 37
rect -35 71 35 109
rect -35 37 -19 71
rect 19 37 35 71
rect -35 21 35 37
rect 93 71 163 109
rect 93 37 109 71
rect 147 37 163 71
rect 93 21 163 37
rect 221 71 291 109
rect 221 37 237 71
rect 275 37 291 71
rect 221 21 291 37
rect 349 71 419 109
rect 349 37 365 71
rect 403 37 419 71
rect 349 21 419 37
rect 477 71 547 109
rect 477 37 493 71
rect 531 37 547 71
rect 477 21 547 37
rect 605 71 675 109
rect 605 37 621 71
rect 659 37 675 71
rect 605 21 675 37
rect 733 71 803 109
rect 733 37 749 71
rect 787 37 803 71
rect 733 21 803 37
rect 861 71 931 109
rect 861 37 877 71
rect 915 37 931 71
rect 861 21 931 37
rect 989 71 1059 109
rect 989 37 1005 71
rect 1043 37 1059 71
rect 989 21 1059 37
rect -1059 -37 -989 -21
rect -1059 -71 -1043 -37
rect -1005 -71 -989 -37
rect -1059 -109 -989 -71
rect -931 -37 -861 -21
rect -931 -71 -915 -37
rect -877 -71 -861 -37
rect -931 -109 -861 -71
rect -803 -37 -733 -21
rect -803 -71 -787 -37
rect -749 -71 -733 -37
rect -803 -109 -733 -71
rect -675 -37 -605 -21
rect -675 -71 -659 -37
rect -621 -71 -605 -37
rect -675 -109 -605 -71
rect -547 -37 -477 -21
rect -547 -71 -531 -37
rect -493 -71 -477 -37
rect -547 -109 -477 -71
rect -419 -37 -349 -21
rect -419 -71 -403 -37
rect -365 -71 -349 -37
rect -419 -109 -349 -71
rect -291 -37 -221 -21
rect -291 -71 -275 -37
rect -237 -71 -221 -37
rect -291 -109 -221 -71
rect -163 -37 -93 -21
rect -163 -71 -147 -37
rect -109 -71 -93 -37
rect -163 -109 -93 -71
rect -35 -37 35 -21
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -35 -109 35 -71
rect 93 -37 163 -21
rect 93 -71 109 -37
rect 147 -71 163 -37
rect 93 -109 163 -71
rect 221 -37 291 -21
rect 221 -71 237 -37
rect 275 -71 291 -37
rect 221 -109 291 -71
rect 349 -37 419 -21
rect 349 -71 365 -37
rect 403 -71 419 -37
rect 349 -109 419 -71
rect 477 -37 547 -21
rect 477 -71 493 -37
rect 531 -71 547 -37
rect 477 -109 547 -71
rect 605 -37 675 -21
rect 605 -71 621 -37
rect 659 -71 675 -37
rect 605 -109 675 -71
rect 733 -37 803 -21
rect 733 -71 749 -37
rect 787 -71 803 -37
rect 733 -109 803 -71
rect 861 -37 931 -21
rect 861 -71 877 -37
rect 915 -71 931 -37
rect 861 -109 931 -71
rect 989 -37 1059 -21
rect 989 -71 1005 -37
rect 1043 -71 1059 -37
rect 989 -109 1059 -71
rect -1059 -647 -989 -609
rect -1059 -681 -1043 -647
rect -1005 -681 -989 -647
rect -1059 -697 -989 -681
rect -931 -647 -861 -609
rect -931 -681 -915 -647
rect -877 -681 -861 -647
rect -931 -697 -861 -681
rect -803 -647 -733 -609
rect -803 -681 -787 -647
rect -749 -681 -733 -647
rect -803 -697 -733 -681
rect -675 -647 -605 -609
rect -675 -681 -659 -647
rect -621 -681 -605 -647
rect -675 -697 -605 -681
rect -547 -647 -477 -609
rect -547 -681 -531 -647
rect -493 -681 -477 -647
rect -547 -697 -477 -681
rect -419 -647 -349 -609
rect -419 -681 -403 -647
rect -365 -681 -349 -647
rect -419 -697 -349 -681
rect -291 -647 -221 -609
rect -291 -681 -275 -647
rect -237 -681 -221 -647
rect -291 -697 -221 -681
rect -163 -647 -93 -609
rect -163 -681 -147 -647
rect -109 -681 -93 -647
rect -163 -697 -93 -681
rect -35 -647 35 -609
rect -35 -681 -19 -647
rect 19 -681 35 -647
rect -35 -697 35 -681
rect 93 -647 163 -609
rect 93 -681 109 -647
rect 147 -681 163 -647
rect 93 -697 163 -681
rect 221 -647 291 -609
rect 221 -681 237 -647
rect 275 -681 291 -647
rect 221 -697 291 -681
rect 349 -647 419 -609
rect 349 -681 365 -647
rect 403 -681 419 -647
rect 349 -697 419 -681
rect 477 -647 547 -609
rect 477 -681 493 -647
rect 531 -681 547 -647
rect 477 -697 547 -681
rect 605 -647 675 -609
rect 605 -681 621 -647
rect 659 -681 675 -647
rect 605 -697 675 -681
rect 733 -647 803 -609
rect 733 -681 749 -647
rect 787 -681 803 -647
rect 733 -697 803 -681
rect 861 -647 931 -609
rect 861 -681 877 -647
rect 915 -681 931 -647
rect 861 -697 931 -681
rect 989 -647 1059 -609
rect 989 -681 1005 -647
rect 1043 -681 1059 -647
rect 989 -697 1059 -681
<< polycont >>
rect -1043 647 -1005 681
rect -915 647 -877 681
rect -787 647 -749 681
rect -659 647 -621 681
rect -531 647 -493 681
rect -403 647 -365 681
rect -275 647 -237 681
rect -147 647 -109 681
rect -19 647 19 681
rect 109 647 147 681
rect 237 647 275 681
rect 365 647 403 681
rect 493 647 531 681
rect 621 647 659 681
rect 749 647 787 681
rect 877 647 915 681
rect 1005 647 1043 681
rect -1043 37 -1005 71
rect -915 37 -877 71
rect -787 37 -749 71
rect -659 37 -621 71
rect -531 37 -493 71
rect -403 37 -365 71
rect -275 37 -237 71
rect -147 37 -109 71
rect -19 37 19 71
rect 109 37 147 71
rect 237 37 275 71
rect 365 37 403 71
rect 493 37 531 71
rect 621 37 659 71
rect 749 37 787 71
rect 877 37 915 71
rect 1005 37 1043 71
rect -1043 -71 -1005 -37
rect -915 -71 -877 -37
rect -787 -71 -749 -37
rect -659 -71 -621 -37
rect -531 -71 -493 -37
rect -403 -71 -365 -37
rect -275 -71 -237 -37
rect -147 -71 -109 -37
rect -19 -71 19 -37
rect 109 -71 147 -37
rect 237 -71 275 -37
rect 365 -71 403 -37
rect 493 -71 531 -37
rect 621 -71 659 -37
rect 749 -71 787 -37
rect 877 -71 915 -37
rect 1005 -71 1043 -37
rect -1043 -681 -1005 -647
rect -915 -681 -877 -647
rect -787 -681 -749 -647
rect -659 -681 -621 -647
rect -531 -681 -493 -647
rect -403 -681 -365 -647
rect -275 -681 -237 -647
rect -147 -681 -109 -647
rect -19 -681 19 -647
rect 109 -681 147 -647
rect 237 -681 275 -647
rect 365 -681 403 -647
rect 493 -681 531 -647
rect 621 -681 659 -647
rect 749 -681 787 -647
rect 877 -681 915 -647
rect 1005 -681 1043 -647
<< locali >>
rect -1219 749 -1123 783
rect 1123 749 1219 783
rect -1219 687 -1185 749
rect 1185 687 1219 749
rect -1059 647 -1043 681
rect -1005 647 -989 681
rect -931 647 -915 681
rect -877 647 -861 681
rect -803 647 -787 681
rect -749 647 -733 681
rect -675 647 -659 681
rect -621 647 -605 681
rect -547 647 -531 681
rect -493 647 -477 681
rect -419 647 -403 681
rect -365 647 -349 681
rect -291 647 -275 681
rect -237 647 -221 681
rect -163 647 -147 681
rect -109 647 -93 681
rect -35 647 -19 681
rect 19 647 35 681
rect 93 647 109 681
rect 147 647 163 681
rect 221 647 237 681
rect 275 647 291 681
rect 349 647 365 681
rect 403 647 419 681
rect 477 647 493 681
rect 531 647 547 681
rect 605 647 621 681
rect 659 647 675 681
rect 733 647 749 681
rect 787 647 803 681
rect 861 647 877 681
rect 915 647 931 681
rect 989 647 1005 681
rect 1043 647 1059 681
rect -1105 597 -1071 613
rect -1105 105 -1071 121
rect -977 597 -943 613
rect -977 105 -943 121
rect -849 597 -815 613
rect -849 105 -815 121
rect -721 597 -687 613
rect -721 105 -687 121
rect -593 597 -559 613
rect -593 105 -559 121
rect -465 597 -431 613
rect -465 105 -431 121
rect -337 597 -303 613
rect -337 105 -303 121
rect -209 597 -175 613
rect -209 105 -175 121
rect -81 597 -47 613
rect -81 105 -47 121
rect 47 597 81 613
rect 47 105 81 121
rect 175 597 209 613
rect 175 105 209 121
rect 303 597 337 613
rect 303 105 337 121
rect 431 597 465 613
rect 431 105 465 121
rect 559 597 593 613
rect 559 105 593 121
rect 687 597 721 613
rect 687 105 721 121
rect 815 597 849 613
rect 815 105 849 121
rect 943 597 977 613
rect 943 105 977 121
rect 1071 597 1105 613
rect 1071 105 1105 121
rect -1059 37 -1043 71
rect -1005 37 -989 71
rect -931 37 -915 71
rect -877 37 -861 71
rect -803 37 -787 71
rect -749 37 -733 71
rect -675 37 -659 71
rect -621 37 -605 71
rect -547 37 -531 71
rect -493 37 -477 71
rect -419 37 -403 71
rect -365 37 -349 71
rect -291 37 -275 71
rect -237 37 -221 71
rect -163 37 -147 71
rect -109 37 -93 71
rect -35 37 -19 71
rect 19 37 35 71
rect 93 37 109 71
rect 147 37 163 71
rect 221 37 237 71
rect 275 37 291 71
rect 349 37 365 71
rect 403 37 419 71
rect 477 37 493 71
rect 531 37 547 71
rect 605 37 621 71
rect 659 37 675 71
rect 733 37 749 71
rect 787 37 803 71
rect 861 37 877 71
rect 915 37 931 71
rect 989 37 1005 71
rect 1043 37 1059 71
rect -1059 -71 -1043 -37
rect -1005 -71 -989 -37
rect -931 -71 -915 -37
rect -877 -71 -861 -37
rect -803 -71 -787 -37
rect -749 -71 -733 -37
rect -675 -71 -659 -37
rect -621 -71 -605 -37
rect -547 -71 -531 -37
rect -493 -71 -477 -37
rect -419 -71 -403 -37
rect -365 -71 -349 -37
rect -291 -71 -275 -37
rect -237 -71 -221 -37
rect -163 -71 -147 -37
rect -109 -71 -93 -37
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect 93 -71 109 -37
rect 147 -71 163 -37
rect 221 -71 237 -37
rect 275 -71 291 -37
rect 349 -71 365 -37
rect 403 -71 419 -37
rect 477 -71 493 -37
rect 531 -71 547 -37
rect 605 -71 621 -37
rect 659 -71 675 -37
rect 733 -71 749 -37
rect 787 -71 803 -37
rect 861 -71 877 -37
rect 915 -71 931 -37
rect 989 -71 1005 -37
rect 1043 -71 1059 -37
rect -1105 -121 -1071 -105
rect -1105 -613 -1071 -597
rect -977 -121 -943 -105
rect -977 -613 -943 -597
rect -849 -121 -815 -105
rect -849 -613 -815 -597
rect -721 -121 -687 -105
rect -721 -613 -687 -597
rect -593 -121 -559 -105
rect -593 -613 -559 -597
rect -465 -121 -431 -105
rect -465 -613 -431 -597
rect -337 -121 -303 -105
rect -337 -613 -303 -597
rect -209 -121 -175 -105
rect -209 -613 -175 -597
rect -81 -121 -47 -105
rect -81 -613 -47 -597
rect 47 -121 81 -105
rect 47 -613 81 -597
rect 175 -121 209 -105
rect 175 -613 209 -597
rect 303 -121 337 -105
rect 303 -613 337 -597
rect 431 -121 465 -105
rect 431 -613 465 -597
rect 559 -121 593 -105
rect 559 -613 593 -597
rect 687 -121 721 -105
rect 687 -613 721 -597
rect 815 -121 849 -105
rect 815 -613 849 -597
rect 943 -121 977 -105
rect 943 -613 977 -597
rect 1071 -121 1105 -105
rect 1071 -613 1105 -597
rect -1059 -681 -1043 -647
rect -1005 -681 -989 -647
rect -931 -681 -915 -647
rect -877 -681 -861 -647
rect -803 -681 -787 -647
rect -749 -681 -733 -647
rect -675 -681 -659 -647
rect -621 -681 -605 -647
rect -547 -681 -531 -647
rect -493 -681 -477 -647
rect -419 -681 -403 -647
rect -365 -681 -349 -647
rect -291 -681 -275 -647
rect -237 -681 -221 -647
rect -163 -681 -147 -647
rect -109 -681 -93 -647
rect -35 -681 -19 -647
rect 19 -681 35 -647
rect 93 -681 109 -647
rect 147 -681 163 -647
rect 221 -681 237 -647
rect 275 -681 291 -647
rect 349 -681 365 -647
rect 403 -681 419 -647
rect 477 -681 493 -647
rect 531 -681 547 -647
rect 605 -681 621 -647
rect 659 -681 675 -647
rect 733 -681 749 -647
rect 787 -681 803 -647
rect 861 -681 877 -647
rect 915 -681 931 -647
rect 989 -681 1005 -647
rect 1043 -681 1059 -647
rect -1219 -749 -1185 -687
rect 1185 -749 1219 -687
rect -1219 -783 -1123 -749
rect 1123 -783 1219 -749
<< viali >>
rect -1043 647 -1005 681
rect -915 647 -877 681
rect -787 647 -749 681
rect -659 647 -621 681
rect -531 647 -493 681
rect -403 647 -365 681
rect -275 647 -237 681
rect -147 647 -109 681
rect -19 647 19 681
rect 109 647 147 681
rect 237 647 275 681
rect 365 647 403 681
rect 493 647 531 681
rect 621 647 659 681
rect 749 647 787 681
rect 877 647 915 681
rect 1005 647 1043 681
rect -1105 121 -1071 597
rect -977 121 -943 597
rect -849 121 -815 597
rect -721 121 -687 597
rect -593 121 -559 597
rect -465 121 -431 597
rect -337 121 -303 597
rect -209 121 -175 597
rect -81 121 -47 597
rect 47 121 81 597
rect 175 121 209 597
rect 303 121 337 597
rect 431 121 465 597
rect 559 121 593 597
rect 687 121 721 597
rect 815 121 849 597
rect 943 121 977 597
rect 1071 121 1105 597
rect -1043 37 -1005 71
rect -915 37 -877 71
rect -787 37 -749 71
rect -659 37 -621 71
rect -531 37 -493 71
rect -403 37 -365 71
rect -275 37 -237 71
rect -147 37 -109 71
rect -19 37 19 71
rect 109 37 147 71
rect 237 37 275 71
rect 365 37 403 71
rect 493 37 531 71
rect 621 37 659 71
rect 749 37 787 71
rect 877 37 915 71
rect 1005 37 1043 71
rect -1043 -71 -1005 -37
rect -915 -71 -877 -37
rect -787 -71 -749 -37
rect -659 -71 -621 -37
rect -531 -71 -493 -37
rect -403 -71 -365 -37
rect -275 -71 -237 -37
rect -147 -71 -109 -37
rect -19 -71 19 -37
rect 109 -71 147 -37
rect 237 -71 275 -37
rect 365 -71 403 -37
rect 493 -71 531 -37
rect 621 -71 659 -37
rect 749 -71 787 -37
rect 877 -71 915 -37
rect 1005 -71 1043 -37
rect -1105 -597 -1071 -121
rect -977 -597 -943 -121
rect -849 -597 -815 -121
rect -721 -597 -687 -121
rect -593 -597 -559 -121
rect -465 -597 -431 -121
rect -337 -597 -303 -121
rect -209 -597 -175 -121
rect -81 -597 -47 -121
rect 47 -597 81 -121
rect 175 -597 209 -121
rect 303 -597 337 -121
rect 431 -597 465 -121
rect 559 -597 593 -121
rect 687 -597 721 -121
rect 815 -597 849 -121
rect 943 -597 977 -121
rect 1071 -597 1105 -121
rect -1043 -681 -1005 -647
rect -915 -681 -877 -647
rect -787 -681 -749 -647
rect -659 -681 -621 -647
rect -531 -681 -493 -647
rect -403 -681 -365 -647
rect -275 -681 -237 -647
rect -147 -681 -109 -647
rect -19 -681 19 -647
rect 109 -681 147 -647
rect 237 -681 275 -647
rect 365 -681 403 -647
rect 493 -681 531 -647
rect 621 -681 659 -647
rect 749 -681 787 -647
rect 877 -681 915 -647
rect 1005 -681 1043 -647
<< metal1 >>
rect -1055 681 -993 687
rect -1055 647 -1043 681
rect -1005 647 -993 681
rect -1055 641 -993 647
rect -927 681 -865 687
rect -927 647 -915 681
rect -877 647 -865 681
rect -927 641 -865 647
rect -799 681 -737 687
rect -799 647 -787 681
rect -749 647 -737 681
rect -799 641 -737 647
rect -671 681 -609 687
rect -671 647 -659 681
rect -621 647 -609 681
rect -671 641 -609 647
rect -543 681 -481 687
rect -543 647 -531 681
rect -493 647 -481 681
rect -543 641 -481 647
rect -415 681 -353 687
rect -415 647 -403 681
rect -365 647 -353 681
rect -415 641 -353 647
rect -287 681 -225 687
rect -287 647 -275 681
rect -237 647 -225 681
rect -287 641 -225 647
rect -159 681 -97 687
rect -159 647 -147 681
rect -109 647 -97 681
rect -159 641 -97 647
rect -31 681 31 687
rect -31 647 -19 681
rect 19 647 31 681
rect -31 641 31 647
rect 97 681 159 687
rect 97 647 109 681
rect 147 647 159 681
rect 97 641 159 647
rect 225 681 287 687
rect 225 647 237 681
rect 275 647 287 681
rect 225 641 287 647
rect 353 681 415 687
rect 353 647 365 681
rect 403 647 415 681
rect 353 641 415 647
rect 481 681 543 687
rect 481 647 493 681
rect 531 647 543 681
rect 481 641 543 647
rect 609 681 671 687
rect 609 647 621 681
rect 659 647 671 681
rect 609 641 671 647
rect 737 681 799 687
rect 737 647 749 681
rect 787 647 799 681
rect 737 641 799 647
rect 865 681 927 687
rect 865 647 877 681
rect 915 647 927 681
rect 865 641 927 647
rect 993 681 1055 687
rect 993 647 1005 681
rect 1043 647 1055 681
rect 993 641 1055 647
rect -1111 597 -1065 609
rect -1111 121 -1105 597
rect -1071 121 -1065 597
rect -1111 109 -1065 121
rect -983 597 -937 609
rect -983 121 -977 597
rect -943 121 -937 597
rect -983 109 -937 121
rect -855 597 -809 609
rect -855 121 -849 597
rect -815 121 -809 597
rect -855 109 -809 121
rect -727 597 -681 609
rect -727 121 -721 597
rect -687 121 -681 597
rect -727 109 -681 121
rect -599 597 -553 609
rect -599 121 -593 597
rect -559 121 -553 597
rect -599 109 -553 121
rect -471 597 -425 609
rect -471 121 -465 597
rect -431 121 -425 597
rect -471 109 -425 121
rect -343 597 -297 609
rect -343 121 -337 597
rect -303 121 -297 597
rect -343 109 -297 121
rect -215 597 -169 609
rect -215 121 -209 597
rect -175 121 -169 597
rect -215 109 -169 121
rect -87 597 -41 609
rect -87 121 -81 597
rect -47 121 -41 597
rect -87 109 -41 121
rect 41 597 87 609
rect 41 121 47 597
rect 81 121 87 597
rect 41 109 87 121
rect 169 597 215 609
rect 169 121 175 597
rect 209 121 215 597
rect 169 109 215 121
rect 297 597 343 609
rect 297 121 303 597
rect 337 121 343 597
rect 297 109 343 121
rect 425 597 471 609
rect 425 121 431 597
rect 465 121 471 597
rect 425 109 471 121
rect 553 597 599 609
rect 553 121 559 597
rect 593 121 599 597
rect 553 109 599 121
rect 681 597 727 609
rect 681 121 687 597
rect 721 121 727 597
rect 681 109 727 121
rect 809 597 855 609
rect 809 121 815 597
rect 849 121 855 597
rect 809 109 855 121
rect 937 597 983 609
rect 937 121 943 597
rect 977 121 983 597
rect 937 109 983 121
rect 1065 597 1111 609
rect 1065 121 1071 597
rect 1105 121 1111 597
rect 1065 109 1111 121
rect -1055 71 -993 77
rect -1055 37 -1043 71
rect -1005 37 -993 71
rect -1055 31 -993 37
rect -927 71 -865 77
rect -927 37 -915 71
rect -877 37 -865 71
rect -927 31 -865 37
rect -799 71 -737 77
rect -799 37 -787 71
rect -749 37 -737 71
rect -799 31 -737 37
rect -671 71 -609 77
rect -671 37 -659 71
rect -621 37 -609 71
rect -671 31 -609 37
rect -543 71 -481 77
rect -543 37 -531 71
rect -493 37 -481 71
rect -543 31 -481 37
rect -415 71 -353 77
rect -415 37 -403 71
rect -365 37 -353 71
rect -415 31 -353 37
rect -287 71 -225 77
rect -287 37 -275 71
rect -237 37 -225 71
rect -287 31 -225 37
rect -159 71 -97 77
rect -159 37 -147 71
rect -109 37 -97 71
rect -159 31 -97 37
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect 97 71 159 77
rect 97 37 109 71
rect 147 37 159 71
rect 97 31 159 37
rect 225 71 287 77
rect 225 37 237 71
rect 275 37 287 71
rect 225 31 287 37
rect 353 71 415 77
rect 353 37 365 71
rect 403 37 415 71
rect 353 31 415 37
rect 481 71 543 77
rect 481 37 493 71
rect 531 37 543 71
rect 481 31 543 37
rect 609 71 671 77
rect 609 37 621 71
rect 659 37 671 71
rect 609 31 671 37
rect 737 71 799 77
rect 737 37 749 71
rect 787 37 799 71
rect 737 31 799 37
rect 865 71 927 77
rect 865 37 877 71
rect 915 37 927 71
rect 865 31 927 37
rect 993 71 1055 77
rect 993 37 1005 71
rect 1043 37 1055 71
rect 993 31 1055 37
rect -1055 -37 -993 -31
rect -1055 -71 -1043 -37
rect -1005 -71 -993 -37
rect -1055 -77 -993 -71
rect -927 -37 -865 -31
rect -927 -71 -915 -37
rect -877 -71 -865 -37
rect -927 -77 -865 -71
rect -799 -37 -737 -31
rect -799 -71 -787 -37
rect -749 -71 -737 -37
rect -799 -77 -737 -71
rect -671 -37 -609 -31
rect -671 -71 -659 -37
rect -621 -71 -609 -37
rect -671 -77 -609 -71
rect -543 -37 -481 -31
rect -543 -71 -531 -37
rect -493 -71 -481 -37
rect -543 -77 -481 -71
rect -415 -37 -353 -31
rect -415 -71 -403 -37
rect -365 -71 -353 -37
rect -415 -77 -353 -71
rect -287 -37 -225 -31
rect -287 -71 -275 -37
rect -237 -71 -225 -37
rect -287 -77 -225 -71
rect -159 -37 -97 -31
rect -159 -71 -147 -37
rect -109 -71 -97 -37
rect -159 -77 -97 -71
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect 97 -37 159 -31
rect 97 -71 109 -37
rect 147 -71 159 -37
rect 97 -77 159 -71
rect 225 -37 287 -31
rect 225 -71 237 -37
rect 275 -71 287 -37
rect 225 -77 287 -71
rect 353 -37 415 -31
rect 353 -71 365 -37
rect 403 -71 415 -37
rect 353 -77 415 -71
rect 481 -37 543 -31
rect 481 -71 493 -37
rect 531 -71 543 -37
rect 481 -77 543 -71
rect 609 -37 671 -31
rect 609 -71 621 -37
rect 659 -71 671 -37
rect 609 -77 671 -71
rect 737 -37 799 -31
rect 737 -71 749 -37
rect 787 -71 799 -37
rect 737 -77 799 -71
rect 865 -37 927 -31
rect 865 -71 877 -37
rect 915 -71 927 -37
rect 865 -77 927 -71
rect 993 -37 1055 -31
rect 993 -71 1005 -37
rect 1043 -71 1055 -37
rect 993 -77 1055 -71
rect -1111 -121 -1065 -109
rect -1111 -597 -1105 -121
rect -1071 -597 -1065 -121
rect -1111 -609 -1065 -597
rect -983 -121 -937 -109
rect -983 -597 -977 -121
rect -943 -597 -937 -121
rect -983 -609 -937 -597
rect -855 -121 -809 -109
rect -855 -597 -849 -121
rect -815 -597 -809 -121
rect -855 -609 -809 -597
rect -727 -121 -681 -109
rect -727 -597 -721 -121
rect -687 -597 -681 -121
rect -727 -609 -681 -597
rect -599 -121 -553 -109
rect -599 -597 -593 -121
rect -559 -597 -553 -121
rect -599 -609 -553 -597
rect -471 -121 -425 -109
rect -471 -597 -465 -121
rect -431 -597 -425 -121
rect -471 -609 -425 -597
rect -343 -121 -297 -109
rect -343 -597 -337 -121
rect -303 -597 -297 -121
rect -343 -609 -297 -597
rect -215 -121 -169 -109
rect -215 -597 -209 -121
rect -175 -597 -169 -121
rect -215 -609 -169 -597
rect -87 -121 -41 -109
rect -87 -597 -81 -121
rect -47 -597 -41 -121
rect -87 -609 -41 -597
rect 41 -121 87 -109
rect 41 -597 47 -121
rect 81 -597 87 -121
rect 41 -609 87 -597
rect 169 -121 215 -109
rect 169 -597 175 -121
rect 209 -597 215 -121
rect 169 -609 215 -597
rect 297 -121 343 -109
rect 297 -597 303 -121
rect 337 -597 343 -121
rect 297 -609 343 -597
rect 425 -121 471 -109
rect 425 -597 431 -121
rect 465 -597 471 -121
rect 425 -609 471 -597
rect 553 -121 599 -109
rect 553 -597 559 -121
rect 593 -597 599 -121
rect 553 -609 599 -597
rect 681 -121 727 -109
rect 681 -597 687 -121
rect 721 -597 727 -121
rect 681 -609 727 -597
rect 809 -121 855 -109
rect 809 -597 815 -121
rect 849 -597 855 -121
rect 809 -609 855 -597
rect 937 -121 983 -109
rect 937 -597 943 -121
rect 977 -597 983 -121
rect 937 -609 983 -597
rect 1065 -121 1111 -109
rect 1065 -597 1071 -121
rect 1105 -597 1111 -121
rect 1065 -609 1111 -597
rect -1055 -647 -993 -641
rect -1055 -681 -1043 -647
rect -1005 -681 -993 -647
rect -1055 -687 -993 -681
rect -927 -647 -865 -641
rect -927 -681 -915 -647
rect -877 -681 -865 -647
rect -927 -687 -865 -681
rect -799 -647 -737 -641
rect -799 -681 -787 -647
rect -749 -681 -737 -647
rect -799 -687 -737 -681
rect -671 -647 -609 -641
rect -671 -681 -659 -647
rect -621 -681 -609 -647
rect -671 -687 -609 -681
rect -543 -647 -481 -641
rect -543 -681 -531 -647
rect -493 -681 -481 -647
rect -543 -687 -481 -681
rect -415 -647 -353 -641
rect -415 -681 -403 -647
rect -365 -681 -353 -647
rect -415 -687 -353 -681
rect -287 -647 -225 -641
rect -287 -681 -275 -647
rect -237 -681 -225 -647
rect -287 -687 -225 -681
rect -159 -647 -97 -641
rect -159 -681 -147 -647
rect -109 -681 -97 -647
rect -159 -687 -97 -681
rect -31 -647 31 -641
rect -31 -681 -19 -647
rect 19 -681 31 -647
rect -31 -687 31 -681
rect 97 -647 159 -641
rect 97 -681 109 -647
rect 147 -681 159 -647
rect 97 -687 159 -681
rect 225 -647 287 -641
rect 225 -681 237 -647
rect 275 -681 287 -647
rect 225 -687 287 -681
rect 353 -647 415 -641
rect 353 -681 365 -647
rect 403 -681 415 -647
rect 353 -687 415 -681
rect 481 -647 543 -641
rect 481 -681 493 -647
rect 531 -681 543 -647
rect 481 -687 543 -681
rect 609 -647 671 -641
rect 609 -681 621 -647
rect 659 -681 671 -647
rect 609 -687 671 -681
rect 737 -647 799 -641
rect 737 -681 749 -647
rect 787 -681 799 -647
rect 737 -687 799 -681
rect 865 -647 927 -641
rect 865 -681 877 -647
rect 915 -681 927 -647
rect 865 -687 927 -681
rect 993 -647 1055 -641
rect 993 -681 1005 -647
rect 1043 -681 1055 -647
rect 993 -687 1055 -681
<< properties >>
string FIXED_BBOX -1202 -766 1202 766
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.5 l 0.35 m 2 nf 17 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
