magic
tech sky130A
magscale 1 2
timestamp 1730410385
<< nwell >>
rect -365 -1219 365 1219
<< pmos >>
rect -169 -1000 -29 1000
rect 29 -1000 169 1000
<< pdiff >>
rect -227 692 -169 1000
rect -227 -692 -215 692
rect -181 -692 -169 692
rect -227 -1000 -169 -692
rect -29 692 29 1000
rect -29 -692 -17 692
rect 17 -692 29 692
rect -29 -1000 29 -692
rect 169 692 227 1000
rect 169 -692 181 692
rect 215 -692 227 692
rect 169 -1000 227 -692
<< pdiffc >>
rect -215 -692 -181 692
rect -17 -692 17 692
rect 181 -692 215 692
<< nsubdiff >>
rect -329 1149 -163 1183
rect 163 1149 329 1183
rect -329 761 -295 1149
rect -329 -1149 -295 -761
rect 295 761 329 1149
rect 295 -1149 329 -761
rect -329 -1183 -163 -1149
rect 163 -1183 329 -1149
<< nsubdiffcont >>
rect -163 1149 163 1183
rect -329 -761 -295 761
rect 295 -761 329 761
rect -163 -1183 163 -1149
<< poly >>
rect -153 1081 -45 1097
rect -153 1064 -137 1081
rect -169 1047 -137 1064
rect -61 1064 -45 1081
rect 45 1081 153 1097
rect 45 1064 61 1081
rect -61 1047 -29 1064
rect -169 1000 -29 1047
rect 29 1047 61 1064
rect 137 1064 153 1081
rect 137 1047 169 1064
rect 29 1000 169 1047
rect -169 -1047 -29 -1000
rect -169 -1064 -137 -1047
rect -153 -1081 -137 -1064
rect -61 -1064 -29 -1047
rect 29 -1047 169 -1000
rect 29 -1064 61 -1047
rect -61 -1081 -45 -1064
rect -153 -1097 -45 -1081
rect 45 -1081 61 -1064
rect 137 -1064 169 -1047
rect 137 -1081 153 -1064
rect 45 -1097 153 -1081
<< polycont >>
rect -137 1047 -61 1081
rect 61 1047 137 1081
rect -137 -1081 -61 -1047
rect 61 -1081 137 -1047
<< locali >>
rect -329 1149 -207 1183
rect 207 1149 329 1183
rect -329 804 -295 1149
rect 295 804 329 1149
rect -215 692 -181 708
rect -215 -708 -181 -692
rect -17 692 17 708
rect -17 -708 17 -692
rect 181 692 215 708
rect 181 -708 215 -692
rect -329 -1149 -295 -804
rect 295 -1149 329 -804
rect -329 -1183 -207 -1149
rect 207 -1183 329 -1149
<< viali >>
rect -207 1149 -163 1183
rect -163 1149 163 1183
rect 163 1149 207 1183
rect -153 1047 -137 1081
rect -137 1047 -61 1081
rect -61 1047 -45 1081
rect 45 1047 61 1081
rect 61 1047 137 1081
rect 137 1047 153 1081
rect -329 761 -295 804
rect -329 -761 -295 761
rect 295 761 329 804
rect -215 -692 -181 692
rect -17 -692 17 692
rect 181 -692 215 692
rect -329 -804 -295 -761
rect 295 -761 329 761
rect 295 -804 329 -761
rect -153 -1081 -137 -1047
rect -137 -1081 -61 -1047
rect -61 -1081 -45 -1047
rect 45 -1081 61 -1047
rect 61 -1081 137 -1047
rect 137 -1081 153 -1047
rect -207 -1183 -163 -1149
rect -163 -1183 163 -1149
rect 163 -1183 207 -1149
<< metal1 >>
rect -219 1183 219 1189
rect -219 1149 -207 1183
rect 207 1149 219 1183
rect -219 1143 219 1149
rect -165 1081 -33 1087
rect -165 1047 -153 1081
rect -45 1047 -33 1081
rect -165 1041 -33 1047
rect 33 1081 165 1087
rect 33 1047 45 1081
rect 153 1047 165 1081
rect 33 1041 165 1047
rect -335 804 -289 816
rect -335 -804 -329 804
rect -295 -804 -289 804
rect 289 804 335 816
rect -221 692 -175 704
rect -221 -692 -215 692
rect -181 -692 -175 692
rect -221 -704 -175 -692
rect -23 692 23 704
rect -23 -692 -17 692
rect 17 -692 23 692
rect -23 -704 23 -692
rect 175 692 221 704
rect 175 -692 181 692
rect 215 -692 221 692
rect 175 -704 221 -692
rect -335 -816 -289 -804
rect 289 -804 295 804
rect 329 -804 335 804
rect 289 -816 335 -804
rect -165 -1047 -33 -1041
rect -165 -1081 -153 -1047
rect -45 -1081 -33 -1047
rect -165 -1087 -33 -1081
rect 33 -1047 165 -1041
rect 33 -1081 45 -1047
rect 153 -1081 165 -1047
rect 33 -1087 165 -1081
rect -219 -1149 219 -1143
rect -219 -1183 -207 -1149
rect 207 -1183 219 -1149
rect -219 -1189 219 -1183
<< properties >>
string FIXED_BBOX -312 -1166 312 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 0.7 m 1 nf 2 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
