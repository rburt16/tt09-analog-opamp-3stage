magic
tech sky130A
magscale 1 2
timestamp 1729530615
<< nwell >>
rect -554 -4573 554 4573
<< pmos >>
rect -358 2354 -158 4354
rect -100 2354 100 4354
rect 158 2354 358 4354
rect -358 118 -158 2118
rect -100 118 100 2118
rect 158 118 358 2118
rect -358 -2118 -158 -118
rect -100 -2118 100 -118
rect 158 -2118 358 -118
rect -358 -4354 -158 -2354
rect -100 -4354 100 -2354
rect 158 -4354 358 -2354
<< pdiff >>
rect -416 4342 -358 4354
rect -416 2366 -404 4342
rect -370 2366 -358 4342
rect -416 2354 -358 2366
rect -158 4342 -100 4354
rect -158 2366 -146 4342
rect -112 2366 -100 4342
rect -158 2354 -100 2366
rect 100 4342 158 4354
rect 100 2366 112 4342
rect 146 2366 158 4342
rect 100 2354 158 2366
rect 358 4342 416 4354
rect 358 2366 370 4342
rect 404 2366 416 4342
rect 358 2354 416 2366
rect -416 2106 -358 2118
rect -416 130 -404 2106
rect -370 130 -358 2106
rect -416 118 -358 130
rect -158 2106 -100 2118
rect -158 130 -146 2106
rect -112 130 -100 2106
rect -158 118 -100 130
rect 100 2106 158 2118
rect 100 130 112 2106
rect 146 130 158 2106
rect 100 118 158 130
rect 358 2106 416 2118
rect 358 130 370 2106
rect 404 130 416 2106
rect 358 118 416 130
rect -416 -130 -358 -118
rect -416 -2106 -404 -130
rect -370 -2106 -358 -130
rect -416 -2118 -358 -2106
rect -158 -130 -100 -118
rect -158 -2106 -146 -130
rect -112 -2106 -100 -130
rect -158 -2118 -100 -2106
rect 100 -130 158 -118
rect 100 -2106 112 -130
rect 146 -2106 158 -130
rect 100 -2118 158 -2106
rect 358 -130 416 -118
rect 358 -2106 370 -130
rect 404 -2106 416 -130
rect 358 -2118 416 -2106
rect -416 -2366 -358 -2354
rect -416 -4342 -404 -2366
rect -370 -4342 -358 -2366
rect -416 -4354 -358 -4342
rect -158 -2366 -100 -2354
rect -158 -4342 -146 -2366
rect -112 -4342 -100 -2366
rect -158 -4354 -100 -4342
rect 100 -2366 158 -2354
rect 100 -4342 112 -2366
rect 146 -4342 158 -2366
rect 100 -4354 158 -4342
rect 358 -2366 416 -2354
rect 358 -4342 370 -2366
rect 404 -4342 416 -2366
rect 358 -4354 416 -4342
<< pdiffc >>
rect -404 2366 -370 4342
rect -146 2366 -112 4342
rect 112 2366 146 4342
rect 370 2366 404 4342
rect -404 130 -370 2106
rect -146 130 -112 2106
rect 112 130 146 2106
rect 370 130 404 2106
rect -404 -2106 -370 -130
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect 370 -2106 404 -130
rect -404 -4342 -370 -2366
rect -146 -4342 -112 -2366
rect 112 -4342 146 -2366
rect 370 -4342 404 -2366
<< nsubdiff >>
rect -518 4503 -422 4537
rect 422 4503 518 4537
rect -518 4441 -484 4503
rect 484 4441 518 4503
rect -518 -4503 -484 -4441
rect 484 -4503 518 -4441
rect -518 -4537 -422 -4503
rect 422 -4537 518 -4503
<< nsubdiffcont >>
rect -422 4503 422 4537
rect -518 -4441 -484 4441
rect 484 -4441 518 4441
rect -422 -4537 422 -4503
<< poly >>
rect -358 4435 -158 4451
rect -358 4401 -342 4435
rect -174 4401 -158 4435
rect -358 4354 -158 4401
rect -100 4435 100 4451
rect -100 4401 -84 4435
rect 84 4401 100 4435
rect -100 4354 100 4401
rect 158 4435 358 4451
rect 158 4401 174 4435
rect 342 4401 358 4435
rect 158 4354 358 4401
rect -358 2307 -158 2354
rect -358 2273 -342 2307
rect -174 2273 -158 2307
rect -358 2257 -158 2273
rect -100 2307 100 2354
rect -100 2273 -84 2307
rect 84 2273 100 2307
rect -100 2257 100 2273
rect 158 2307 358 2354
rect 158 2273 174 2307
rect 342 2273 358 2307
rect 158 2257 358 2273
rect -358 2199 -158 2215
rect -358 2165 -342 2199
rect -174 2165 -158 2199
rect -358 2118 -158 2165
rect -100 2199 100 2215
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -100 2118 100 2165
rect 158 2199 358 2215
rect 158 2165 174 2199
rect 342 2165 358 2199
rect 158 2118 358 2165
rect -358 71 -158 118
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -118 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -118 358 -71
rect -358 -2165 -158 -2118
rect -358 -2199 -342 -2165
rect -174 -2199 -158 -2165
rect -358 -2215 -158 -2199
rect -100 -2165 100 -2118
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -100 -2215 100 -2199
rect 158 -2165 358 -2118
rect 158 -2199 174 -2165
rect 342 -2199 358 -2165
rect 158 -2215 358 -2199
rect -358 -2273 -158 -2257
rect -358 -2307 -342 -2273
rect -174 -2307 -158 -2273
rect -358 -2354 -158 -2307
rect -100 -2273 100 -2257
rect -100 -2307 -84 -2273
rect 84 -2307 100 -2273
rect -100 -2354 100 -2307
rect 158 -2273 358 -2257
rect 158 -2307 174 -2273
rect 342 -2307 358 -2273
rect 158 -2354 358 -2307
rect -358 -4401 -158 -4354
rect -358 -4435 -342 -4401
rect -174 -4435 -158 -4401
rect -358 -4451 -158 -4435
rect -100 -4401 100 -4354
rect -100 -4435 -84 -4401
rect 84 -4435 100 -4401
rect -100 -4451 100 -4435
rect 158 -4401 358 -4354
rect 158 -4435 174 -4401
rect 342 -4435 358 -4401
rect 158 -4451 358 -4435
<< polycont >>
rect -342 4401 -174 4435
rect -84 4401 84 4435
rect 174 4401 342 4435
rect -342 2273 -174 2307
rect -84 2273 84 2307
rect 174 2273 342 2307
rect -342 2165 -174 2199
rect -84 2165 84 2199
rect 174 2165 342 2199
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect -342 -2199 -174 -2165
rect -84 -2199 84 -2165
rect 174 -2199 342 -2165
rect -342 -2307 -174 -2273
rect -84 -2307 84 -2273
rect 174 -2307 342 -2273
rect -342 -4435 -174 -4401
rect -84 -4435 84 -4401
rect 174 -4435 342 -4401
<< locali >>
rect -518 4503 -422 4537
rect 422 4503 518 4537
rect -518 4441 -484 4503
rect 484 4441 518 4503
rect -358 4401 -342 4435
rect -174 4401 -158 4435
rect -100 4401 -84 4435
rect 84 4401 100 4435
rect 158 4401 174 4435
rect 342 4401 358 4435
rect -404 4342 -370 4358
rect -404 2350 -370 2366
rect -146 4342 -112 4358
rect -146 2350 -112 2366
rect 112 4342 146 4358
rect 112 2350 146 2366
rect 370 4342 404 4358
rect 370 2350 404 2366
rect -358 2273 -342 2307
rect -174 2273 -158 2307
rect -100 2273 -84 2307
rect 84 2273 100 2307
rect 158 2273 174 2307
rect 342 2273 358 2307
rect -358 2165 -342 2199
rect -174 2165 -158 2199
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect 158 2165 174 2199
rect 342 2165 358 2199
rect -404 2106 -370 2122
rect -404 114 -370 130
rect -146 2106 -112 2122
rect -146 114 -112 130
rect 112 2106 146 2122
rect 112 114 146 130
rect 370 2106 404 2122
rect 370 114 404 130
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect -404 -130 -370 -114
rect -404 -2122 -370 -2106
rect -146 -130 -112 -114
rect -146 -2122 -112 -2106
rect 112 -130 146 -114
rect 112 -2122 146 -2106
rect 370 -130 404 -114
rect 370 -2122 404 -2106
rect -358 -2199 -342 -2165
rect -174 -2199 -158 -2165
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect 158 -2199 174 -2165
rect 342 -2199 358 -2165
rect -358 -2307 -342 -2273
rect -174 -2307 -158 -2273
rect -100 -2307 -84 -2273
rect 84 -2307 100 -2273
rect 158 -2307 174 -2273
rect 342 -2307 358 -2273
rect -404 -2366 -370 -2350
rect -404 -4358 -370 -4342
rect -146 -2366 -112 -2350
rect -146 -4358 -112 -4342
rect 112 -2366 146 -2350
rect 112 -4358 146 -4342
rect 370 -2366 404 -2350
rect 370 -4358 404 -4342
rect -358 -4435 -342 -4401
rect -174 -4435 -158 -4401
rect -100 -4435 -84 -4401
rect 84 -4435 100 -4401
rect 158 -4435 174 -4401
rect 342 -4435 358 -4401
rect -518 -4503 -484 -4441
rect 484 -4503 518 -4441
rect -518 -4537 -422 -4503
rect 422 -4537 518 -4503
<< viali >>
rect -342 4401 -174 4435
rect -84 4401 84 4435
rect 174 4401 342 4435
rect -404 2366 -370 4342
rect -146 2366 -112 4342
rect 112 2366 146 4342
rect 370 2366 404 4342
rect -342 2273 -174 2307
rect -84 2273 84 2307
rect 174 2273 342 2307
rect -342 2165 -174 2199
rect -84 2165 84 2199
rect 174 2165 342 2199
rect -404 130 -370 2106
rect -146 130 -112 2106
rect 112 130 146 2106
rect 370 130 404 2106
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect -404 -2106 -370 -130
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect 370 -2106 404 -130
rect -342 -2199 -174 -2165
rect -84 -2199 84 -2165
rect 174 -2199 342 -2165
rect -342 -2307 -174 -2273
rect -84 -2307 84 -2273
rect 174 -2307 342 -2273
rect -404 -4342 -370 -2366
rect -146 -4342 -112 -2366
rect 112 -4342 146 -2366
rect 370 -4342 404 -2366
rect -342 -4435 -174 -4401
rect -84 -4435 84 -4401
rect 174 -4435 342 -4401
<< metal1 >>
rect -354 4435 -162 4441
rect -354 4401 -342 4435
rect -174 4401 -162 4435
rect -354 4395 -162 4401
rect -96 4435 96 4441
rect -96 4401 -84 4435
rect 84 4401 96 4435
rect -96 4395 96 4401
rect 162 4435 354 4441
rect 162 4401 174 4435
rect 342 4401 354 4435
rect 162 4395 354 4401
rect -410 4342 -364 4354
rect -410 2366 -404 4342
rect -370 2366 -364 4342
rect -410 2354 -364 2366
rect -152 4342 -106 4354
rect -152 2366 -146 4342
rect -112 2366 -106 4342
rect -152 2354 -106 2366
rect 106 4342 152 4354
rect 106 2366 112 4342
rect 146 2366 152 4342
rect 106 2354 152 2366
rect 364 4342 410 4354
rect 364 2366 370 4342
rect 404 2366 410 4342
rect 364 2354 410 2366
rect -354 2307 -162 2313
rect -354 2273 -342 2307
rect -174 2273 -162 2307
rect -354 2267 -162 2273
rect -96 2307 96 2313
rect -96 2273 -84 2307
rect 84 2273 96 2307
rect -96 2267 96 2273
rect 162 2307 354 2313
rect 162 2273 174 2307
rect 342 2273 354 2307
rect 162 2267 354 2273
rect -354 2199 -162 2205
rect -354 2165 -342 2199
rect -174 2165 -162 2199
rect -354 2159 -162 2165
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect 162 2199 354 2205
rect 162 2165 174 2199
rect 342 2165 354 2199
rect 162 2159 354 2165
rect -410 2106 -364 2118
rect -410 130 -404 2106
rect -370 130 -364 2106
rect -410 118 -364 130
rect -152 2106 -106 2118
rect -152 130 -146 2106
rect -112 130 -106 2106
rect -152 118 -106 130
rect 106 2106 152 2118
rect 106 130 112 2106
rect 146 130 152 2106
rect 106 118 152 130
rect 364 2106 410 2118
rect 364 130 370 2106
rect 404 130 410 2106
rect 364 118 410 130
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect -410 -130 -364 -118
rect -410 -2106 -404 -130
rect -370 -2106 -364 -130
rect -410 -2118 -364 -2106
rect -152 -130 -106 -118
rect -152 -2106 -146 -130
rect -112 -2106 -106 -130
rect -152 -2118 -106 -2106
rect 106 -130 152 -118
rect 106 -2106 112 -130
rect 146 -2106 152 -130
rect 106 -2118 152 -2106
rect 364 -130 410 -118
rect 364 -2106 370 -130
rect 404 -2106 410 -130
rect 364 -2118 410 -2106
rect -354 -2165 -162 -2159
rect -354 -2199 -342 -2165
rect -174 -2199 -162 -2165
rect -354 -2205 -162 -2199
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
rect 162 -2165 354 -2159
rect 162 -2199 174 -2165
rect 342 -2199 354 -2165
rect 162 -2205 354 -2199
rect -354 -2273 -162 -2267
rect -354 -2307 -342 -2273
rect -174 -2307 -162 -2273
rect -354 -2313 -162 -2307
rect -96 -2273 96 -2267
rect -96 -2307 -84 -2273
rect 84 -2307 96 -2273
rect -96 -2313 96 -2307
rect 162 -2273 354 -2267
rect 162 -2307 174 -2273
rect 342 -2307 354 -2273
rect 162 -2313 354 -2307
rect -410 -2366 -364 -2354
rect -410 -4342 -404 -2366
rect -370 -4342 -364 -2366
rect -410 -4354 -364 -4342
rect -152 -2366 -106 -2354
rect -152 -4342 -146 -2366
rect -112 -4342 -106 -2366
rect -152 -4354 -106 -4342
rect 106 -2366 152 -2354
rect 106 -4342 112 -2366
rect 146 -4342 152 -2366
rect 106 -4354 152 -4342
rect 364 -2366 410 -2354
rect 364 -4342 370 -2366
rect 404 -4342 410 -2366
rect 364 -4354 410 -4342
rect -354 -4401 -162 -4395
rect -354 -4435 -342 -4401
rect -174 -4435 -162 -4401
rect -354 -4441 -162 -4435
rect -96 -4401 96 -4395
rect -96 -4435 -84 -4401
rect 84 -4435 96 -4401
rect -96 -4441 96 -4435
rect 162 -4401 354 -4395
rect 162 -4435 174 -4401
rect 342 -4435 354 -4401
rect 162 -4441 354 -4435
<< properties >>
string FIXED_BBOX -501 -4520 501 4520
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 4 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
