magic
tech sky130A
magscale 1 2
timestamp 1729267537
<< pwell >>
rect -596 -1919 596 1919
<< nmoslvt >>
rect -400 109 400 1709
rect -400 -1709 400 -109
<< ndiff >>
rect -458 1697 -400 1709
rect -458 121 -446 1697
rect -412 121 -400 1697
rect -458 109 -400 121
rect 400 1697 458 1709
rect 400 121 412 1697
rect 446 121 458 1697
rect 400 109 458 121
rect -458 -121 -400 -109
rect -458 -1697 -446 -121
rect -412 -1697 -400 -121
rect -458 -1709 -400 -1697
rect 400 -121 458 -109
rect 400 -1697 412 -121
rect 446 -1697 458 -121
rect 400 -1709 458 -1697
<< ndiffc >>
rect -446 121 -412 1697
rect 412 121 446 1697
rect -446 -1697 -412 -121
rect 412 -1697 446 -121
<< psubdiff >>
rect -560 1849 -464 1883
rect 464 1849 560 1883
rect -560 1787 -526 1849
rect 526 1787 560 1849
rect -560 -1849 -526 -1787
rect 526 -1849 560 -1787
rect -560 -1883 -464 -1849
rect 464 -1883 560 -1849
<< psubdiffcont >>
rect -464 1849 464 1883
rect -560 -1787 -526 1787
rect 526 -1787 560 1787
rect -464 -1883 464 -1849
<< poly >>
rect -400 1781 400 1797
rect -400 1747 -384 1781
rect 384 1747 400 1781
rect -400 1709 400 1747
rect -400 71 400 109
rect -400 37 -384 71
rect 384 37 400 71
rect -400 21 400 37
rect -400 -37 400 -21
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -400 -109 400 -71
rect -400 -1747 400 -1709
rect -400 -1781 -384 -1747
rect 384 -1781 400 -1747
rect -400 -1797 400 -1781
<< polycont >>
rect -384 1747 384 1781
rect -384 37 384 71
rect -384 -71 384 -37
rect -384 -1781 384 -1747
<< locali >>
rect -560 1849 -464 1883
rect 464 1849 560 1883
rect -560 1787 -526 1849
rect 526 1787 560 1849
rect -400 1747 -384 1781
rect 384 1747 400 1781
rect -446 1697 -412 1713
rect -446 105 -412 121
rect 412 1697 446 1713
rect 412 105 446 121
rect -400 37 -384 71
rect 384 37 400 71
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -446 -121 -412 -105
rect -446 -1713 -412 -1697
rect 412 -121 446 -105
rect 412 -1713 446 -1697
rect -400 -1781 -384 -1747
rect 384 -1781 400 -1747
rect -560 -1849 -526 -1787
rect 526 -1849 560 -1787
rect -560 -1883 -464 -1849
rect 464 -1883 560 -1849
<< viali >>
rect -384 1747 384 1781
rect -446 121 -412 1697
rect 412 121 446 1697
rect -384 37 384 71
rect -384 -71 384 -37
rect -446 -1697 -412 -121
rect 412 -1697 446 -121
rect -384 -1781 384 -1747
<< metal1 >>
rect -396 1781 396 1787
rect -396 1747 -384 1781
rect 384 1747 396 1781
rect -396 1741 396 1747
rect -452 1697 -406 1709
rect -452 121 -446 1697
rect -412 121 -406 1697
rect -452 109 -406 121
rect 406 1697 452 1709
rect 406 121 412 1697
rect 446 121 452 1697
rect 406 109 452 121
rect -396 71 396 77
rect -396 37 -384 71
rect 384 37 396 71
rect -396 31 396 37
rect -396 -37 396 -31
rect -396 -71 -384 -37
rect 384 -71 396 -37
rect -396 -77 396 -71
rect -452 -121 -406 -109
rect -452 -1697 -446 -121
rect -412 -1697 -406 -121
rect -452 -1709 -406 -1697
rect 406 -121 452 -109
rect 406 -1697 412 -121
rect 446 -1697 452 -121
rect 406 -1709 452 -1697
rect -396 -1747 396 -1741
rect -396 -1781 -384 -1747
rect 384 -1781 396 -1747
rect -396 -1787 396 -1781
<< properties >>
string FIXED_BBOX -543 -1866 543 1866
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8.0 l 4.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
