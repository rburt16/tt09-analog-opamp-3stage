magic
tech sky130A
magscale 1 2
timestamp 1728061155
<< metal3 >>
rect -13104 2712 -6732 2740
rect -13104 -2712 -6816 2712
rect -6752 -2712 -6732 2712
rect -13104 -2740 -6732 -2712
rect -6492 2712 -120 2740
rect -6492 -2712 -204 2712
rect -140 -2712 -120 2712
rect -6492 -2740 -120 -2712
rect 120 2712 6492 2740
rect 120 -2712 6408 2712
rect 6472 -2712 6492 2712
rect 120 -2740 6492 -2712
rect 6732 2712 13104 2740
rect 6732 -2712 13020 2712
rect 13084 -2712 13104 2712
rect 6732 -2740 13104 -2712
<< via3 >>
rect -6816 -2712 -6752 2712
rect -204 -2712 -140 2712
rect 6408 -2712 6472 2712
rect 13020 -2712 13084 2712
<< mimcap >>
rect -13064 2660 -7064 2700
rect -13064 -2660 -13024 2660
rect -7104 -2660 -7064 2660
rect -13064 -2700 -7064 -2660
rect -6452 2660 -452 2700
rect -6452 -2660 -6412 2660
rect -492 -2660 -452 2660
rect -6452 -2700 -452 -2660
rect 160 2660 6160 2700
rect 160 -2660 200 2660
rect 6120 -2660 6160 2660
rect 160 -2700 6160 -2660
rect 6772 2660 12772 2700
rect 6772 -2660 6812 2660
rect 12732 -2660 12772 2660
rect 6772 -2700 12772 -2660
<< mimcapcontact >>
rect -13024 -2660 -7104 2660
rect -6412 -2660 -492 2660
rect 200 -2660 6120 2660
rect 6812 -2660 12732 2660
<< metal4 >>
rect -6832 2712 -6736 2728
rect -13025 2660 -7103 2661
rect -13025 -2660 -13024 2660
rect -7104 -2660 -7103 2660
rect -13025 -2661 -7103 -2660
rect -6832 -2712 -6816 2712
rect -6752 -2712 -6736 2712
rect -220 2712 -124 2728
rect -6413 2660 -491 2661
rect -6413 -2660 -6412 2660
rect -492 -2660 -491 2660
rect -6413 -2661 -491 -2660
rect -6832 -2728 -6736 -2712
rect -220 -2712 -204 2712
rect -140 -2712 -124 2712
rect 6392 2712 6488 2728
rect 199 2660 6121 2661
rect 199 -2660 200 2660
rect 6120 -2660 6121 2660
rect 199 -2661 6121 -2660
rect -220 -2728 -124 -2712
rect 6392 -2712 6408 2712
rect 6472 -2712 6488 2712
rect 13004 2712 13100 2728
rect 6811 2660 12733 2661
rect 6811 -2660 6812 2660
rect 12732 -2660 12733 2660
rect 6811 -2661 12733 -2660
rect 6392 -2728 6488 -2712
rect 13004 -2712 13020 2712
rect 13084 -2712 13100 2712
rect 13004 -2728 13100 -2712
<< properties >>
string FIXED_BBOX 6732 -2740 12812 2740
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 27.0 val 1.641k carea 2.00 cperi 0.19 nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
