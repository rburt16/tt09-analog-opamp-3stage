magic
tech sky130A
magscale 1 2
timestamp 1730139296
<< error_p >>
rect -671 2199 -609 2205
rect -543 2199 -481 2205
rect -415 2199 -353 2205
rect -287 2199 -225 2205
rect -159 2199 -97 2205
rect -31 2199 31 2205
rect 97 2199 159 2205
rect 225 2199 287 2205
rect 353 2199 415 2205
rect 481 2199 543 2205
rect 609 2199 671 2205
rect -671 2165 -659 2199
rect -543 2165 -531 2199
rect -415 2165 -403 2199
rect -287 2165 -275 2199
rect -159 2165 -147 2199
rect -31 2165 -19 2199
rect 97 2165 109 2199
rect 225 2165 237 2199
rect 353 2165 365 2199
rect 481 2165 493 2199
rect 609 2165 621 2199
rect -671 2159 -609 2165
rect -543 2159 -481 2165
rect -415 2159 -353 2165
rect -287 2159 -225 2165
rect -159 2159 -97 2165
rect -31 2159 31 2165
rect 97 2159 159 2165
rect 225 2159 287 2165
rect 353 2159 415 2165
rect 481 2159 543 2165
rect 609 2159 671 2165
rect -671 71 -609 77
rect -543 71 -481 77
rect -415 71 -353 77
rect -287 71 -225 77
rect -159 71 -97 77
rect -31 71 31 77
rect 97 71 159 77
rect 225 71 287 77
rect 353 71 415 77
rect 481 71 543 77
rect 609 71 671 77
rect -671 37 -659 71
rect -543 37 -531 71
rect -415 37 -403 71
rect -287 37 -275 71
rect -159 37 -147 71
rect -31 37 -19 71
rect 97 37 109 71
rect 225 37 237 71
rect 353 37 365 71
rect 481 37 493 71
rect 609 37 621 71
rect -671 31 -609 37
rect -543 31 -481 37
rect -415 31 -353 37
rect -287 31 -225 37
rect -159 31 -97 37
rect -31 31 31 37
rect 97 31 159 37
rect 225 31 287 37
rect 353 31 415 37
rect 481 31 543 37
rect 609 31 671 37
rect -671 -37 -609 -31
rect -543 -37 -481 -31
rect -415 -37 -353 -31
rect -287 -37 -225 -31
rect -159 -37 -97 -31
rect -31 -37 31 -31
rect 97 -37 159 -31
rect 225 -37 287 -31
rect 353 -37 415 -31
rect 481 -37 543 -31
rect 609 -37 671 -31
rect -671 -71 -659 -37
rect -543 -71 -531 -37
rect -415 -71 -403 -37
rect -287 -71 -275 -37
rect -159 -71 -147 -37
rect -31 -71 -19 -37
rect 97 -71 109 -37
rect 225 -71 237 -37
rect 353 -71 365 -37
rect 481 -71 493 -37
rect 609 -71 621 -37
rect -671 -77 -609 -71
rect -543 -77 -481 -71
rect -415 -77 -353 -71
rect -287 -77 -225 -71
rect -159 -77 -97 -71
rect -31 -77 31 -71
rect 97 -77 159 -71
rect 225 -77 287 -71
rect 353 -77 415 -71
rect 481 -77 543 -71
rect 609 -77 671 -71
rect -671 -2165 -609 -2159
rect -543 -2165 -481 -2159
rect -415 -2165 -353 -2159
rect -287 -2165 -225 -2159
rect -159 -2165 -97 -2159
rect -31 -2165 31 -2159
rect 97 -2165 159 -2159
rect 225 -2165 287 -2159
rect 353 -2165 415 -2159
rect 481 -2165 543 -2159
rect 609 -2165 671 -2159
rect -671 -2199 -659 -2165
rect -543 -2199 -531 -2165
rect -415 -2199 -403 -2165
rect -287 -2199 -275 -2165
rect -159 -2199 -147 -2165
rect -31 -2199 -19 -2165
rect 97 -2199 109 -2165
rect 225 -2199 237 -2165
rect 353 -2199 365 -2165
rect 481 -2199 493 -2165
rect 609 -2199 621 -2165
rect -671 -2205 -609 -2199
rect -543 -2205 -481 -2199
rect -415 -2205 -353 -2199
rect -287 -2205 -225 -2199
rect -159 -2205 -97 -2199
rect -31 -2205 31 -2199
rect 97 -2205 159 -2199
rect 225 -2205 287 -2199
rect 353 -2205 415 -2199
rect 481 -2205 543 -2199
rect 609 -2205 671 -2199
<< nwell >>
rect -871 -2337 871 2337
<< pmoslvt >>
rect -675 118 -605 2118
rect -547 118 -477 2118
rect -419 118 -349 2118
rect -291 118 -221 2118
rect -163 118 -93 2118
rect -35 118 35 2118
rect 93 118 163 2118
rect 221 118 291 2118
rect 349 118 419 2118
rect 477 118 547 2118
rect 605 118 675 2118
rect -675 -2118 -605 -118
rect -547 -2118 -477 -118
rect -419 -2118 -349 -118
rect -291 -2118 -221 -118
rect -163 -2118 -93 -118
rect -35 -2118 35 -118
rect 93 -2118 163 -118
rect 221 -2118 291 -118
rect 349 -2118 419 -118
rect 477 -2118 547 -118
rect 605 -2118 675 -118
<< pdiff >>
rect -733 1810 -675 2118
rect -733 426 -721 1810
rect -687 426 -675 1810
rect -733 118 -675 426
rect -605 1810 -547 2118
rect -605 426 -593 1810
rect -559 426 -547 1810
rect -605 118 -547 426
rect -477 1810 -419 2118
rect -477 426 -465 1810
rect -431 426 -419 1810
rect -477 118 -419 426
rect -349 1810 -291 2118
rect -349 426 -337 1810
rect -303 426 -291 1810
rect -349 118 -291 426
rect -221 1810 -163 2118
rect -221 426 -209 1810
rect -175 426 -163 1810
rect -221 118 -163 426
rect -93 1810 -35 2118
rect -93 426 -81 1810
rect -47 426 -35 1810
rect -93 118 -35 426
rect 35 1810 93 2118
rect 35 426 47 1810
rect 81 426 93 1810
rect 35 118 93 426
rect 163 1810 221 2118
rect 163 426 175 1810
rect 209 426 221 1810
rect 163 118 221 426
rect 291 1810 349 2118
rect 291 426 303 1810
rect 337 426 349 1810
rect 291 118 349 426
rect 419 1810 477 2118
rect 419 426 431 1810
rect 465 426 477 1810
rect 419 118 477 426
rect 547 1810 605 2118
rect 547 426 559 1810
rect 593 426 605 1810
rect 547 118 605 426
rect 675 1810 733 2118
rect 675 426 687 1810
rect 721 426 733 1810
rect 675 118 733 426
rect -733 -426 -675 -118
rect -733 -1810 -721 -426
rect -687 -1810 -675 -426
rect -733 -2118 -675 -1810
rect -605 -426 -547 -118
rect -605 -1810 -593 -426
rect -559 -1810 -547 -426
rect -605 -2118 -547 -1810
rect -477 -426 -419 -118
rect -477 -1810 -465 -426
rect -431 -1810 -419 -426
rect -477 -2118 -419 -1810
rect -349 -426 -291 -118
rect -349 -1810 -337 -426
rect -303 -1810 -291 -426
rect -349 -2118 -291 -1810
rect -221 -426 -163 -118
rect -221 -1810 -209 -426
rect -175 -1810 -163 -426
rect -221 -2118 -163 -1810
rect -93 -426 -35 -118
rect -93 -1810 -81 -426
rect -47 -1810 -35 -426
rect -93 -2118 -35 -1810
rect 35 -426 93 -118
rect 35 -1810 47 -426
rect 81 -1810 93 -426
rect 35 -2118 93 -1810
rect 163 -426 221 -118
rect 163 -1810 175 -426
rect 209 -1810 221 -426
rect 163 -2118 221 -1810
rect 291 -426 349 -118
rect 291 -1810 303 -426
rect 337 -1810 349 -426
rect 291 -2118 349 -1810
rect 419 -426 477 -118
rect 419 -1810 431 -426
rect 465 -1810 477 -426
rect 419 -2118 477 -1810
rect 547 -426 605 -118
rect 547 -1810 559 -426
rect 593 -1810 605 -426
rect 547 -2118 605 -1810
rect 675 -426 733 -118
rect 675 -1810 687 -426
rect 721 -1810 733 -426
rect 675 -2118 733 -1810
<< pdiffc >>
rect -721 426 -687 1810
rect -593 426 -559 1810
rect -465 426 -431 1810
rect -337 426 -303 1810
rect -209 426 -175 1810
rect -81 426 -47 1810
rect 47 426 81 1810
rect 175 426 209 1810
rect 303 426 337 1810
rect 431 426 465 1810
rect 559 426 593 1810
rect 687 426 721 1810
rect -721 -1810 -687 -426
rect -593 -1810 -559 -426
rect -465 -1810 -431 -426
rect -337 -1810 -303 -426
rect -209 -1810 -175 -426
rect -81 -1810 -47 -426
rect 47 -1810 81 -426
rect 175 -1810 209 -426
rect 303 -1810 337 -426
rect 431 -1810 465 -426
rect 559 -1810 593 -426
rect 687 -1810 721 -426
<< nsubdiff >>
rect -835 2267 835 2301
rect -835 1544 -801 2267
rect -835 -2267 -801 -1544
rect 801 -2267 835 2267
rect -835 -2301 835 -2267
<< nsubdiffcont >>
rect -835 -1544 -801 1544
<< poly >>
rect -673 2199 -607 2215
rect -673 2182 -657 2199
rect -675 2165 -657 2182
rect -623 2182 -607 2199
rect -545 2199 -479 2215
rect -545 2182 -529 2199
rect -623 2165 -605 2182
rect -675 2118 -605 2165
rect -547 2165 -529 2182
rect -495 2182 -479 2199
rect -417 2199 -351 2215
rect -417 2182 -401 2199
rect -495 2165 -477 2182
rect -547 2118 -477 2165
rect -419 2165 -401 2182
rect -367 2182 -351 2199
rect -289 2199 -223 2215
rect -289 2182 -273 2199
rect -367 2165 -349 2182
rect -419 2118 -349 2165
rect -291 2165 -273 2182
rect -239 2182 -223 2199
rect -161 2199 -95 2215
rect -161 2182 -145 2199
rect -239 2165 -221 2182
rect -291 2118 -221 2165
rect -163 2165 -145 2182
rect -111 2182 -95 2199
rect -33 2199 33 2215
rect -33 2182 -17 2199
rect -111 2165 -93 2182
rect -163 2118 -93 2165
rect -35 2165 -17 2182
rect 17 2182 33 2199
rect 95 2199 161 2215
rect 95 2182 111 2199
rect 17 2165 35 2182
rect -35 2118 35 2165
rect 93 2165 111 2182
rect 145 2182 161 2199
rect 223 2199 289 2215
rect 223 2182 239 2199
rect 145 2165 163 2182
rect 93 2118 163 2165
rect 221 2165 239 2182
rect 273 2182 289 2199
rect 351 2199 417 2215
rect 351 2182 367 2199
rect 273 2165 291 2182
rect 221 2118 291 2165
rect 349 2165 367 2182
rect 401 2182 417 2199
rect 479 2199 545 2215
rect 479 2182 495 2199
rect 401 2165 419 2182
rect 349 2118 419 2165
rect 477 2165 495 2182
rect 529 2182 545 2199
rect 607 2199 673 2215
rect 607 2182 623 2199
rect 529 2165 547 2182
rect 477 2118 547 2165
rect 605 2165 623 2182
rect 657 2182 673 2199
rect 657 2165 675 2182
rect 605 2118 675 2165
rect -675 71 -605 118
rect -675 54 -657 71
rect -673 37 -657 54
rect -623 54 -605 71
rect -547 71 -477 118
rect -547 54 -529 71
rect -623 37 -607 54
rect -673 21 -607 37
rect -545 37 -529 54
rect -495 54 -477 71
rect -419 71 -349 118
rect -419 54 -401 71
rect -495 37 -479 54
rect -545 21 -479 37
rect -417 37 -401 54
rect -367 54 -349 71
rect -291 71 -221 118
rect -291 54 -273 71
rect -367 37 -351 54
rect -417 21 -351 37
rect -289 37 -273 54
rect -239 54 -221 71
rect -163 71 -93 118
rect -163 54 -145 71
rect -239 37 -223 54
rect -289 21 -223 37
rect -161 37 -145 54
rect -111 54 -93 71
rect -35 71 35 118
rect -35 54 -17 71
rect -111 37 -95 54
rect -161 21 -95 37
rect -33 37 -17 54
rect 17 54 35 71
rect 93 71 163 118
rect 93 54 111 71
rect 17 37 33 54
rect -33 21 33 37
rect 95 37 111 54
rect 145 54 163 71
rect 221 71 291 118
rect 221 54 239 71
rect 145 37 161 54
rect 95 21 161 37
rect 223 37 239 54
rect 273 54 291 71
rect 349 71 419 118
rect 349 54 367 71
rect 273 37 289 54
rect 223 21 289 37
rect 351 37 367 54
rect 401 54 419 71
rect 477 71 547 118
rect 477 54 495 71
rect 401 37 417 54
rect 351 21 417 37
rect 479 37 495 54
rect 529 54 547 71
rect 605 71 675 118
rect 605 54 623 71
rect 529 37 545 54
rect 479 21 545 37
rect 607 37 623 54
rect 657 54 675 71
rect 657 37 673 54
rect 607 21 673 37
rect -673 -37 -607 -21
rect -673 -54 -657 -37
rect -675 -71 -657 -54
rect -623 -54 -607 -37
rect -545 -37 -479 -21
rect -545 -54 -529 -37
rect -623 -71 -605 -54
rect -675 -118 -605 -71
rect -547 -71 -529 -54
rect -495 -54 -479 -37
rect -417 -37 -351 -21
rect -417 -54 -401 -37
rect -495 -71 -477 -54
rect -547 -118 -477 -71
rect -419 -71 -401 -54
rect -367 -54 -351 -37
rect -289 -37 -223 -21
rect -289 -54 -273 -37
rect -367 -71 -349 -54
rect -419 -118 -349 -71
rect -291 -71 -273 -54
rect -239 -54 -223 -37
rect -161 -37 -95 -21
rect -161 -54 -145 -37
rect -239 -71 -221 -54
rect -291 -118 -221 -71
rect -163 -71 -145 -54
rect -111 -54 -95 -37
rect -33 -37 33 -21
rect -33 -54 -17 -37
rect -111 -71 -93 -54
rect -163 -118 -93 -71
rect -35 -71 -17 -54
rect 17 -54 33 -37
rect 95 -37 161 -21
rect 95 -54 111 -37
rect 17 -71 35 -54
rect -35 -118 35 -71
rect 93 -71 111 -54
rect 145 -54 161 -37
rect 223 -37 289 -21
rect 223 -54 239 -37
rect 145 -71 163 -54
rect 93 -118 163 -71
rect 221 -71 239 -54
rect 273 -54 289 -37
rect 351 -37 417 -21
rect 351 -54 367 -37
rect 273 -71 291 -54
rect 221 -118 291 -71
rect 349 -71 367 -54
rect 401 -54 417 -37
rect 479 -37 545 -21
rect 479 -54 495 -37
rect 401 -71 419 -54
rect 349 -118 419 -71
rect 477 -71 495 -54
rect 529 -54 545 -37
rect 607 -37 673 -21
rect 607 -54 623 -37
rect 529 -71 547 -54
rect 477 -118 547 -71
rect 605 -71 623 -54
rect 657 -54 673 -37
rect 657 -71 675 -54
rect 605 -118 675 -71
rect -675 -2165 -605 -2118
rect -675 -2182 -657 -2165
rect -673 -2199 -657 -2182
rect -623 -2182 -605 -2165
rect -547 -2165 -477 -2118
rect -547 -2182 -529 -2165
rect -623 -2199 -607 -2182
rect -673 -2215 -607 -2199
rect -545 -2199 -529 -2182
rect -495 -2182 -477 -2165
rect -419 -2165 -349 -2118
rect -419 -2182 -401 -2165
rect -495 -2199 -479 -2182
rect -545 -2215 -479 -2199
rect -417 -2199 -401 -2182
rect -367 -2182 -349 -2165
rect -291 -2165 -221 -2118
rect -291 -2182 -273 -2165
rect -367 -2199 -351 -2182
rect -417 -2215 -351 -2199
rect -289 -2199 -273 -2182
rect -239 -2182 -221 -2165
rect -163 -2165 -93 -2118
rect -163 -2182 -145 -2165
rect -239 -2199 -223 -2182
rect -289 -2215 -223 -2199
rect -161 -2199 -145 -2182
rect -111 -2182 -93 -2165
rect -35 -2165 35 -2118
rect -35 -2182 -17 -2165
rect -111 -2199 -95 -2182
rect -161 -2215 -95 -2199
rect -33 -2199 -17 -2182
rect 17 -2182 35 -2165
rect 93 -2165 163 -2118
rect 93 -2182 111 -2165
rect 17 -2199 33 -2182
rect -33 -2215 33 -2199
rect 95 -2199 111 -2182
rect 145 -2182 163 -2165
rect 221 -2165 291 -2118
rect 221 -2182 239 -2165
rect 145 -2199 161 -2182
rect 95 -2215 161 -2199
rect 223 -2199 239 -2182
rect 273 -2182 291 -2165
rect 349 -2165 419 -2118
rect 349 -2182 367 -2165
rect 273 -2199 289 -2182
rect 223 -2215 289 -2199
rect 351 -2199 367 -2182
rect 401 -2182 419 -2165
rect 477 -2165 547 -2118
rect 477 -2182 495 -2165
rect 401 -2199 417 -2182
rect 351 -2215 417 -2199
rect 479 -2199 495 -2182
rect 529 -2182 547 -2165
rect 605 -2165 675 -2118
rect 605 -2182 623 -2165
rect 529 -2199 545 -2182
rect 479 -2215 545 -2199
rect 607 -2199 623 -2182
rect 657 -2182 675 -2165
rect 657 -2199 673 -2182
rect 607 -2215 673 -2199
<< polycont >>
rect -657 2165 -623 2199
rect -529 2165 -495 2199
rect -401 2165 -367 2199
rect -273 2165 -239 2199
rect -145 2165 -111 2199
rect -17 2165 17 2199
rect 111 2165 145 2199
rect 239 2165 273 2199
rect 367 2165 401 2199
rect 495 2165 529 2199
rect 623 2165 657 2199
rect -657 37 -623 71
rect -529 37 -495 71
rect -401 37 -367 71
rect -273 37 -239 71
rect -145 37 -111 71
rect -17 37 17 71
rect 111 37 145 71
rect 239 37 273 71
rect 367 37 401 71
rect 495 37 529 71
rect 623 37 657 71
rect -657 -71 -623 -37
rect -529 -71 -495 -37
rect -401 -71 -367 -37
rect -273 -71 -239 -37
rect -145 -71 -111 -37
rect -17 -71 17 -37
rect 111 -71 145 -37
rect 239 -71 273 -37
rect 367 -71 401 -37
rect 495 -71 529 -37
rect 623 -71 657 -37
rect -657 -2199 -623 -2165
rect -529 -2199 -495 -2165
rect -401 -2199 -367 -2165
rect -273 -2199 -239 -2165
rect -145 -2199 -111 -2165
rect -17 -2199 17 -2165
rect 111 -2199 145 -2165
rect 239 -2199 273 -2165
rect 367 -2199 401 -2165
rect 495 -2199 529 -2165
rect 623 -2199 657 -2165
<< locali >>
rect -835 2267 835 2301
rect -835 1587 -801 2267
rect -673 2165 -659 2199
rect -621 2165 -607 2199
rect -545 2165 -531 2199
rect -493 2165 -479 2199
rect -417 2165 -403 2199
rect -365 2165 -351 2199
rect -289 2165 -275 2199
rect -237 2165 -223 2199
rect -161 2165 -147 2199
rect -109 2165 -95 2199
rect -33 2165 -19 2199
rect 19 2165 33 2199
rect 95 2165 109 2199
rect 147 2165 161 2199
rect 223 2165 237 2199
rect 275 2165 289 2199
rect 351 2165 365 2199
rect 403 2165 417 2199
rect 479 2165 493 2199
rect 531 2165 545 2199
rect 607 2165 621 2199
rect 659 2165 673 2199
rect -721 1810 -687 1826
rect -721 410 -687 426
rect -593 1810 -559 1826
rect -593 410 -559 426
rect -465 1810 -431 1826
rect -465 410 -431 426
rect -337 1810 -303 1826
rect -337 410 -303 426
rect -209 1810 -175 1826
rect -209 410 -175 426
rect -81 1810 -47 1826
rect -81 410 -47 426
rect 47 1810 81 1826
rect 47 410 81 426
rect 175 1810 209 1826
rect 175 410 209 426
rect 303 1810 337 1826
rect 303 410 337 426
rect 431 1810 465 1826
rect 431 410 465 426
rect 559 1810 593 1826
rect 559 410 593 426
rect 687 1810 721 1826
rect 687 410 721 426
rect -673 37 -659 71
rect -621 37 -607 71
rect -545 37 -531 71
rect -493 37 -479 71
rect -417 37 -403 71
rect -365 37 -351 71
rect -289 37 -275 71
rect -237 37 -223 71
rect -161 37 -147 71
rect -109 37 -95 71
rect -33 37 -19 71
rect 19 37 33 71
rect 95 37 109 71
rect 147 37 161 71
rect 223 37 237 71
rect 275 37 289 71
rect 351 37 365 71
rect 403 37 417 71
rect 479 37 493 71
rect 531 37 545 71
rect 607 37 621 71
rect 659 37 673 71
rect -673 -71 -659 -37
rect -621 -71 -607 -37
rect -545 -71 -531 -37
rect -493 -71 -479 -37
rect -417 -71 -403 -37
rect -365 -71 -351 -37
rect -289 -71 -275 -37
rect -237 -71 -223 -37
rect -161 -71 -147 -37
rect -109 -71 -95 -37
rect -33 -71 -19 -37
rect 19 -71 33 -37
rect 95 -71 109 -37
rect 147 -71 161 -37
rect 223 -71 237 -37
rect 275 -71 289 -37
rect 351 -71 365 -37
rect 403 -71 417 -37
rect 479 -71 493 -37
rect 531 -71 545 -37
rect 607 -71 621 -37
rect 659 -71 673 -37
rect -835 -2267 -801 -1587
rect -721 -426 -687 -410
rect -721 -1826 -687 -1810
rect -593 -426 -559 -410
rect -593 -1826 -559 -1810
rect -465 -426 -431 -410
rect -465 -1826 -431 -1810
rect -337 -426 -303 -410
rect -337 -1826 -303 -1810
rect -209 -426 -175 -410
rect -209 -1826 -175 -1810
rect -81 -426 -47 -410
rect -81 -1826 -47 -1810
rect 47 -426 81 -410
rect 47 -1826 81 -1810
rect 175 -426 209 -410
rect 175 -1826 209 -1810
rect 303 -426 337 -410
rect 303 -1826 337 -1810
rect 431 -426 465 -410
rect 431 -1826 465 -1810
rect 559 -426 593 -410
rect 559 -1826 593 -1810
rect 687 -426 721 -410
rect 687 -1826 721 -1810
rect -673 -2199 -659 -2165
rect -621 -2199 -607 -2165
rect -545 -2199 -531 -2165
rect -493 -2199 -479 -2165
rect -417 -2199 -403 -2165
rect -365 -2199 -351 -2165
rect -289 -2199 -275 -2165
rect -237 -2199 -223 -2165
rect -161 -2199 -147 -2165
rect -109 -2199 -95 -2165
rect -33 -2199 -19 -2165
rect 19 -2199 33 -2165
rect 95 -2199 109 -2165
rect 147 -2199 161 -2165
rect 223 -2199 237 -2165
rect 275 -2199 289 -2165
rect 351 -2199 365 -2165
rect 403 -2199 417 -2165
rect 479 -2199 493 -2165
rect 531 -2199 545 -2165
rect 607 -2199 621 -2165
rect 659 -2199 673 -2165
rect 801 -2267 835 2267
rect -835 -2301 835 -2267
<< viali >>
rect -659 2165 -657 2199
rect -657 2165 -623 2199
rect -623 2165 -621 2199
rect -531 2165 -529 2199
rect -529 2165 -495 2199
rect -495 2165 -493 2199
rect -403 2165 -401 2199
rect -401 2165 -367 2199
rect -367 2165 -365 2199
rect -275 2165 -273 2199
rect -273 2165 -239 2199
rect -239 2165 -237 2199
rect -147 2165 -145 2199
rect -145 2165 -111 2199
rect -111 2165 -109 2199
rect -19 2165 -17 2199
rect -17 2165 17 2199
rect 17 2165 19 2199
rect 109 2165 111 2199
rect 111 2165 145 2199
rect 145 2165 147 2199
rect 237 2165 239 2199
rect 239 2165 273 2199
rect 273 2165 275 2199
rect 365 2165 367 2199
rect 367 2165 401 2199
rect 401 2165 403 2199
rect 493 2165 495 2199
rect 495 2165 529 2199
rect 529 2165 531 2199
rect 621 2165 623 2199
rect 623 2165 657 2199
rect 657 2165 659 2199
rect -835 1544 -801 1587
rect -835 -1544 -801 1544
rect -721 426 -687 1810
rect -593 426 -559 1810
rect -465 426 -431 1810
rect -337 426 -303 1810
rect -209 426 -175 1810
rect -81 426 -47 1810
rect 47 426 81 1810
rect 175 426 209 1810
rect 303 426 337 1810
rect 431 426 465 1810
rect 559 426 593 1810
rect 687 426 721 1810
rect -659 37 -657 71
rect -657 37 -623 71
rect -623 37 -621 71
rect -531 37 -529 71
rect -529 37 -495 71
rect -495 37 -493 71
rect -403 37 -401 71
rect -401 37 -367 71
rect -367 37 -365 71
rect -275 37 -273 71
rect -273 37 -239 71
rect -239 37 -237 71
rect -147 37 -145 71
rect -145 37 -111 71
rect -111 37 -109 71
rect -19 37 -17 71
rect -17 37 17 71
rect 17 37 19 71
rect 109 37 111 71
rect 111 37 145 71
rect 145 37 147 71
rect 237 37 239 71
rect 239 37 273 71
rect 273 37 275 71
rect 365 37 367 71
rect 367 37 401 71
rect 401 37 403 71
rect 493 37 495 71
rect 495 37 529 71
rect 529 37 531 71
rect 621 37 623 71
rect 623 37 657 71
rect 657 37 659 71
rect -659 -71 -657 -37
rect -657 -71 -623 -37
rect -623 -71 -621 -37
rect -531 -71 -529 -37
rect -529 -71 -495 -37
rect -495 -71 -493 -37
rect -403 -71 -401 -37
rect -401 -71 -367 -37
rect -367 -71 -365 -37
rect -275 -71 -273 -37
rect -273 -71 -239 -37
rect -239 -71 -237 -37
rect -147 -71 -145 -37
rect -145 -71 -111 -37
rect -111 -71 -109 -37
rect -19 -71 -17 -37
rect -17 -71 17 -37
rect 17 -71 19 -37
rect 109 -71 111 -37
rect 111 -71 145 -37
rect 145 -71 147 -37
rect 237 -71 239 -37
rect 239 -71 273 -37
rect 273 -71 275 -37
rect 365 -71 367 -37
rect 367 -71 401 -37
rect 401 -71 403 -37
rect 493 -71 495 -37
rect 495 -71 529 -37
rect 529 -71 531 -37
rect 621 -71 623 -37
rect 623 -71 657 -37
rect 657 -71 659 -37
rect -835 -1587 -801 -1544
rect -721 -1810 -687 -426
rect -593 -1810 -559 -426
rect -465 -1810 -431 -426
rect -337 -1810 -303 -426
rect -209 -1810 -175 -426
rect -81 -1810 -47 -426
rect 47 -1810 81 -426
rect 175 -1810 209 -426
rect 303 -1810 337 -426
rect 431 -1810 465 -426
rect 559 -1810 593 -426
rect 687 -1810 721 -426
rect -659 -2199 -657 -2165
rect -657 -2199 -623 -2165
rect -623 -2199 -621 -2165
rect -531 -2199 -529 -2165
rect -529 -2199 -495 -2165
rect -495 -2199 -493 -2165
rect -403 -2199 -401 -2165
rect -401 -2199 -367 -2165
rect -367 -2199 -365 -2165
rect -275 -2199 -273 -2165
rect -273 -2199 -239 -2165
rect -239 -2199 -237 -2165
rect -147 -2199 -145 -2165
rect -145 -2199 -111 -2165
rect -111 -2199 -109 -2165
rect -19 -2199 -17 -2165
rect -17 -2199 17 -2165
rect 17 -2199 19 -2165
rect 109 -2199 111 -2165
rect 111 -2199 145 -2165
rect 145 -2199 147 -2165
rect 237 -2199 239 -2165
rect 239 -2199 273 -2165
rect 273 -2199 275 -2165
rect 365 -2199 367 -2165
rect 367 -2199 401 -2165
rect 401 -2199 403 -2165
rect 493 -2199 495 -2165
rect 495 -2199 529 -2165
rect 529 -2199 531 -2165
rect 621 -2199 623 -2165
rect 623 -2199 657 -2165
rect 657 -2199 659 -2165
<< metal1 >>
rect -671 2199 -609 2205
rect -671 2165 -659 2199
rect -621 2165 -609 2199
rect -671 2159 -609 2165
rect -543 2199 -481 2205
rect -543 2165 -531 2199
rect -493 2165 -481 2199
rect -543 2159 -481 2165
rect -415 2199 -353 2205
rect -415 2165 -403 2199
rect -365 2165 -353 2199
rect -415 2159 -353 2165
rect -287 2199 -225 2205
rect -287 2165 -275 2199
rect -237 2165 -225 2199
rect -287 2159 -225 2165
rect -159 2199 -97 2205
rect -159 2165 -147 2199
rect -109 2165 -97 2199
rect -159 2159 -97 2165
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect 19 2165 31 2199
rect -31 2159 31 2165
rect 97 2199 159 2205
rect 97 2165 109 2199
rect 147 2165 159 2199
rect 97 2159 159 2165
rect 225 2199 287 2205
rect 225 2165 237 2199
rect 275 2165 287 2199
rect 225 2159 287 2165
rect 353 2199 415 2205
rect 353 2165 365 2199
rect 403 2165 415 2199
rect 353 2159 415 2165
rect 481 2199 543 2205
rect 481 2165 493 2199
rect 531 2165 543 2199
rect 481 2159 543 2165
rect 609 2199 671 2205
rect 609 2165 621 2199
rect 659 2165 671 2199
rect 609 2159 671 2165
rect -727 1810 -681 1822
rect -841 1587 -795 1599
rect -841 -1587 -835 1587
rect -801 -1587 -795 1587
rect -727 426 -721 1810
rect -687 426 -681 1810
rect -727 414 -681 426
rect -599 1810 -553 1822
rect -599 426 -593 1810
rect -559 426 -553 1810
rect -599 414 -553 426
rect -471 1810 -425 1822
rect -471 426 -465 1810
rect -431 426 -425 1810
rect -471 414 -425 426
rect -343 1810 -297 1822
rect -343 426 -337 1810
rect -303 426 -297 1810
rect -343 414 -297 426
rect -215 1810 -169 1822
rect -215 426 -209 1810
rect -175 426 -169 1810
rect -215 414 -169 426
rect -87 1810 -41 1822
rect -87 426 -81 1810
rect -47 426 -41 1810
rect -87 414 -41 426
rect 41 1810 87 1822
rect 41 426 47 1810
rect 81 426 87 1810
rect 41 414 87 426
rect 169 1810 215 1822
rect 169 426 175 1810
rect 209 426 215 1810
rect 169 414 215 426
rect 297 1810 343 1822
rect 297 426 303 1810
rect 337 426 343 1810
rect 297 414 343 426
rect 425 1810 471 1822
rect 425 426 431 1810
rect 465 426 471 1810
rect 425 414 471 426
rect 553 1810 599 1822
rect 553 426 559 1810
rect 593 426 599 1810
rect 553 414 599 426
rect 681 1810 727 1822
rect 681 426 687 1810
rect 721 426 727 1810
rect 681 414 727 426
rect -671 71 -609 77
rect -671 37 -659 71
rect -621 37 -609 71
rect -671 31 -609 37
rect -543 71 -481 77
rect -543 37 -531 71
rect -493 37 -481 71
rect -543 31 -481 37
rect -415 71 -353 77
rect -415 37 -403 71
rect -365 37 -353 71
rect -415 31 -353 37
rect -287 71 -225 77
rect -287 37 -275 71
rect -237 37 -225 71
rect -287 31 -225 37
rect -159 71 -97 77
rect -159 37 -147 71
rect -109 37 -97 71
rect -159 31 -97 37
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect 97 71 159 77
rect 97 37 109 71
rect 147 37 159 71
rect 97 31 159 37
rect 225 71 287 77
rect 225 37 237 71
rect 275 37 287 71
rect 225 31 287 37
rect 353 71 415 77
rect 353 37 365 71
rect 403 37 415 71
rect 353 31 415 37
rect 481 71 543 77
rect 481 37 493 71
rect 531 37 543 71
rect 481 31 543 37
rect 609 71 671 77
rect 609 37 621 71
rect 659 37 671 71
rect 609 31 671 37
rect -671 -37 -609 -31
rect -671 -71 -659 -37
rect -621 -71 -609 -37
rect -671 -77 -609 -71
rect -543 -37 -481 -31
rect -543 -71 -531 -37
rect -493 -71 -481 -37
rect -543 -77 -481 -71
rect -415 -37 -353 -31
rect -415 -71 -403 -37
rect -365 -71 -353 -37
rect -415 -77 -353 -71
rect -287 -37 -225 -31
rect -287 -71 -275 -37
rect -237 -71 -225 -37
rect -287 -77 -225 -71
rect -159 -37 -97 -31
rect -159 -71 -147 -37
rect -109 -71 -97 -37
rect -159 -77 -97 -71
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect 97 -37 159 -31
rect 97 -71 109 -37
rect 147 -71 159 -37
rect 97 -77 159 -71
rect 225 -37 287 -31
rect 225 -71 237 -37
rect 275 -71 287 -37
rect 225 -77 287 -71
rect 353 -37 415 -31
rect 353 -71 365 -37
rect 403 -71 415 -37
rect 353 -77 415 -71
rect 481 -37 543 -31
rect 481 -71 493 -37
rect 531 -71 543 -37
rect 481 -77 543 -71
rect 609 -37 671 -31
rect 609 -71 621 -37
rect 659 -71 671 -37
rect 609 -77 671 -71
rect -841 -1599 -795 -1587
rect -727 -426 -681 -414
rect -727 -1810 -721 -426
rect -687 -1810 -681 -426
rect -727 -1822 -681 -1810
rect -599 -426 -553 -414
rect -599 -1810 -593 -426
rect -559 -1810 -553 -426
rect -599 -1822 -553 -1810
rect -471 -426 -425 -414
rect -471 -1810 -465 -426
rect -431 -1810 -425 -426
rect -471 -1822 -425 -1810
rect -343 -426 -297 -414
rect -343 -1810 -337 -426
rect -303 -1810 -297 -426
rect -343 -1822 -297 -1810
rect -215 -426 -169 -414
rect -215 -1810 -209 -426
rect -175 -1810 -169 -426
rect -215 -1822 -169 -1810
rect -87 -426 -41 -414
rect -87 -1810 -81 -426
rect -47 -1810 -41 -426
rect -87 -1822 -41 -1810
rect 41 -426 87 -414
rect 41 -1810 47 -426
rect 81 -1810 87 -426
rect 41 -1822 87 -1810
rect 169 -426 215 -414
rect 169 -1810 175 -426
rect 209 -1810 215 -426
rect 169 -1822 215 -1810
rect 297 -426 343 -414
rect 297 -1810 303 -426
rect 337 -1810 343 -426
rect 297 -1822 343 -1810
rect 425 -426 471 -414
rect 425 -1810 431 -426
rect 465 -1810 471 -426
rect 425 -1822 471 -1810
rect 553 -426 599 -414
rect 553 -1810 559 -426
rect 593 -1810 599 -426
rect 553 -1822 599 -1810
rect 681 -426 727 -414
rect 681 -1810 687 -426
rect 721 -1810 727 -426
rect 681 -1822 727 -1810
rect -671 -2165 -609 -2159
rect -671 -2199 -659 -2165
rect -621 -2199 -609 -2165
rect -671 -2205 -609 -2199
rect -543 -2165 -481 -2159
rect -543 -2199 -531 -2165
rect -493 -2199 -481 -2165
rect -543 -2205 -481 -2199
rect -415 -2165 -353 -2159
rect -415 -2199 -403 -2165
rect -365 -2199 -353 -2165
rect -415 -2205 -353 -2199
rect -287 -2165 -225 -2159
rect -287 -2199 -275 -2165
rect -237 -2199 -225 -2165
rect -287 -2205 -225 -2199
rect -159 -2165 -97 -2159
rect -159 -2199 -147 -2165
rect -109 -2199 -97 -2165
rect -159 -2205 -97 -2199
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect 19 -2199 31 -2165
rect -31 -2205 31 -2199
rect 97 -2165 159 -2159
rect 97 -2199 109 -2165
rect 147 -2199 159 -2165
rect 97 -2205 159 -2199
rect 225 -2165 287 -2159
rect 225 -2199 237 -2165
rect 275 -2199 287 -2165
rect 225 -2205 287 -2199
rect 353 -2165 415 -2159
rect 353 -2199 365 -2165
rect 403 -2199 415 -2165
rect 353 -2205 415 -2199
rect 481 -2165 543 -2159
rect 481 -2199 493 -2165
rect 531 -2199 543 -2165
rect 481 -2205 543 -2199
rect 609 -2165 671 -2159
rect 609 -2199 621 -2165
rect 659 -2199 671 -2165
rect 609 -2205 671 -2199
<< properties >>
string FIXED_BBOX -818 -2284 818 2284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 2 nf 11 diffcov 70 polycov 70 guard 1 glc 1 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 0 viagr 0 viagl 70 viagt 0
<< end >>
