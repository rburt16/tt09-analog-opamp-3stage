magic
tech sky130A
magscale 1 2
timestamp 1729267537
<< nwell >>
rect -365 -1219 365 1219
<< pmos >>
rect -169 -1000 -29 1000
rect 29 -1000 169 1000
<< pdiff >>
rect -227 988 -169 1000
rect -227 -988 -215 988
rect -181 -988 -169 988
rect -227 -1000 -169 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 169 988 227 1000
rect 169 -988 181 988
rect 215 -988 227 988
rect 169 -1000 227 -988
<< pdiffc >>
rect -215 -988 -181 988
rect -17 -988 17 988
rect 181 -988 215 988
<< nsubdiff >>
rect -329 1149 -233 1183
rect 233 1149 329 1183
rect -329 1087 -295 1149
rect 295 1087 329 1149
rect -329 -1149 -295 -1087
rect 295 -1149 329 -1087
rect -329 -1183 -233 -1149
rect 233 -1183 329 -1149
<< nsubdiffcont >>
rect -233 1149 233 1183
rect -329 -1087 -295 1087
rect 295 -1087 329 1087
rect -233 -1183 233 -1149
<< poly >>
rect -169 1081 -29 1097
rect -169 1047 -153 1081
rect -45 1047 -29 1081
rect -169 1000 -29 1047
rect 29 1081 169 1097
rect 29 1047 45 1081
rect 153 1047 169 1081
rect 29 1000 169 1047
rect -169 -1047 -29 -1000
rect -169 -1081 -153 -1047
rect -45 -1081 -29 -1047
rect -169 -1097 -29 -1081
rect 29 -1047 169 -1000
rect 29 -1081 45 -1047
rect 153 -1081 169 -1047
rect 29 -1097 169 -1081
<< polycont >>
rect -153 1047 -45 1081
rect 45 1047 153 1081
rect -153 -1081 -45 -1047
rect 45 -1081 153 -1047
<< locali >>
rect -329 1149 -233 1183
rect 233 1149 329 1183
rect -329 1087 -295 1149
rect 295 1087 329 1149
rect -169 1047 -153 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 153 1047 169 1081
rect -215 988 -181 1004
rect -215 -1004 -181 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 181 988 215 1004
rect 181 -1004 215 -988
rect -169 -1081 -153 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 153 -1081 169 -1047
rect -329 -1149 -295 -1087
rect 295 -1149 329 -1087
rect -329 -1183 -233 -1149
rect 233 -1183 329 -1149
<< viali >>
rect -153 1047 -45 1081
rect 45 1047 153 1081
rect -215 -988 -181 988
rect -17 -988 17 988
rect 181 -988 215 988
rect -153 -1081 -45 -1047
rect 45 -1081 153 -1047
<< metal1 >>
rect -165 1081 -33 1087
rect -165 1047 -153 1081
rect -45 1047 -33 1081
rect -165 1041 -33 1047
rect 33 1081 165 1087
rect 33 1047 45 1081
rect 153 1047 165 1081
rect 33 1041 165 1047
rect -221 988 -175 1000
rect -221 -988 -215 988
rect -181 -988 -175 988
rect -221 -1000 -175 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 175 988 221 1000
rect 175 -988 181 988
rect 215 -988 221 988
rect 175 -1000 221 -988
rect -165 -1047 -33 -1041
rect -165 -1081 -153 -1047
rect -45 -1081 -33 -1047
rect -165 -1087 -33 -1081
rect 33 -1047 165 -1041
rect 33 -1081 45 -1047
rect 153 -1081 165 -1047
rect 33 -1087 165 -1081
<< properties >>
string FIXED_BBOX -312 -1166 312 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 0.7 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
