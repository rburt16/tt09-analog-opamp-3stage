magic
tech sky130A
timestamp 1728938857
<< pwell >>
rect -298 -255 298 255
<< nmoslvt >>
rect -200 -150 200 150
<< ndiff >>
rect -229 144 -200 150
rect -229 -144 -223 144
rect -206 -144 -200 144
rect -229 -150 -200 -144
rect 200 144 229 150
rect 200 -144 206 144
rect 223 -144 229 144
rect 200 -150 229 -144
<< ndiffc >>
rect -223 -144 -206 144
rect 206 -144 223 144
<< psubdiff >>
rect -280 220 -232 237
rect 232 220 280 237
rect -280 189 -263 220
rect 263 189 280 220
rect -280 -220 -263 -189
rect 263 -220 280 -189
rect -280 -237 -232 -220
rect 232 -237 280 -220
<< psubdiffcont >>
rect -232 220 232 237
rect -280 -189 -263 189
rect 263 -189 280 189
rect -232 -237 232 -220
<< poly >>
rect -200 186 200 194
rect -200 169 -192 186
rect 192 169 200 186
rect -200 150 200 169
rect -200 -169 200 -150
rect -200 -186 -192 -169
rect 192 -186 200 -169
rect -200 -194 200 -186
<< polycont >>
rect -192 169 192 186
rect -192 -186 192 -169
<< locali >>
rect -280 220 -232 237
rect 232 220 280 237
rect -280 189 -263 220
rect 263 189 280 220
rect -200 169 -192 186
rect 192 169 200 186
rect -223 144 -206 152
rect -223 -152 -206 -144
rect 206 144 223 152
rect 206 -152 223 -144
rect -200 -186 -192 -169
rect 192 -186 200 -169
rect -280 -220 -263 -189
rect 263 -220 280 -189
rect -280 -237 -232 -220
rect 232 -237 280 -220
<< viali >>
rect -192 169 192 186
rect -223 -144 -206 144
rect 206 -144 223 144
rect -192 -186 192 -169
<< metal1 >>
rect -198 186 198 189
rect -198 169 -192 186
rect 192 169 198 186
rect -198 166 198 169
rect -226 144 -203 150
rect -226 -144 -223 144
rect -206 -144 -203 144
rect -226 -150 -203 -144
rect 203 144 226 150
rect 203 -144 206 144
rect 223 -144 226 144
rect 203 -150 226 -144
rect -198 -169 198 -166
rect -198 -186 -192 -169
rect 192 -186 198 -169
rect -198 -189 198 -186
<< properties >>
string FIXED_BBOX -271 -228 271 228
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3.0 l 4.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
