magic
tech sky130A
magscale 1 2
timestamp 1729617920
<< nwell >>
rect -554 -2337 554 2337
<< pmos >>
rect -358 118 -158 2118
rect -100 118 100 2118
rect 158 118 358 2118
rect -358 -2118 -158 -118
rect -100 -2118 100 -118
rect 158 -2118 358 -118
<< pdiff >>
rect -416 2106 -358 2118
rect -416 130 -404 2106
rect -370 130 -358 2106
rect -416 118 -358 130
rect -158 2106 -100 2118
rect -158 130 -146 2106
rect -112 130 -100 2106
rect -158 118 -100 130
rect 100 2106 158 2118
rect 100 130 112 2106
rect 146 130 158 2106
rect 100 118 158 130
rect 358 2106 416 2118
rect 358 130 370 2106
rect 404 130 416 2106
rect 358 118 416 130
rect -416 -130 -358 -118
rect -416 -2106 -404 -130
rect -370 -2106 -358 -130
rect -416 -2118 -358 -2106
rect -158 -130 -100 -118
rect -158 -2106 -146 -130
rect -112 -2106 -100 -130
rect -158 -2118 -100 -2106
rect 100 -130 158 -118
rect 100 -2106 112 -130
rect 146 -2106 158 -130
rect 100 -2118 158 -2106
rect 358 -130 416 -118
rect 358 -2106 370 -130
rect 404 -2106 416 -130
rect 358 -2118 416 -2106
<< pdiffc >>
rect -404 130 -370 2106
rect -146 130 -112 2106
rect 112 130 146 2106
rect 370 130 404 2106
rect -404 -2106 -370 -130
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect 370 -2106 404 -130
<< nsubdiff >>
rect -518 2267 -422 2301
rect 422 2267 518 2301
rect -518 2205 -484 2267
rect 484 2205 518 2267
rect -518 -2267 -484 -2205
rect 484 -2267 518 -2205
rect -518 -2301 -422 -2267
rect 422 -2301 518 -2267
<< nsubdiffcont >>
rect -422 2267 422 2301
rect -518 -2205 -484 2205
rect 484 -2205 518 2205
rect -422 -2301 422 -2267
<< poly >>
rect -358 2199 -158 2215
rect -358 2165 -342 2199
rect -174 2165 -158 2199
rect -358 2118 -158 2165
rect -100 2199 100 2215
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect -100 2118 100 2165
rect 158 2199 358 2215
rect 158 2165 174 2199
rect 342 2165 358 2199
rect 158 2118 358 2165
rect -358 71 -158 118
rect -358 37 -342 71
rect -174 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 174 71
rect 342 37 358 71
rect 158 21 358 37
rect -358 -37 -158 -21
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -358 -118 -158 -71
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect 158 -37 358 -21
rect 158 -71 174 -37
rect 342 -71 358 -37
rect 158 -118 358 -71
rect -358 -2165 -158 -2118
rect -358 -2199 -342 -2165
rect -174 -2199 -158 -2165
rect -358 -2215 -158 -2199
rect -100 -2165 100 -2118
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect -100 -2215 100 -2199
rect 158 -2165 358 -2118
rect 158 -2199 174 -2165
rect 342 -2199 358 -2165
rect 158 -2215 358 -2199
<< polycont >>
rect -342 2165 -174 2199
rect -84 2165 84 2199
rect 174 2165 342 2199
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect -342 -2199 -174 -2165
rect -84 -2199 84 -2165
rect 174 -2199 342 -2165
<< locali >>
rect -518 2267 -422 2301
rect 422 2267 518 2301
rect -518 2205 -484 2267
rect 484 2205 518 2267
rect -358 2165 -342 2199
rect -174 2165 -158 2199
rect -100 2165 -84 2199
rect 84 2165 100 2199
rect 158 2165 174 2199
rect 342 2165 358 2199
rect -404 2106 -370 2122
rect -404 114 -370 130
rect -146 2106 -112 2122
rect -146 114 -112 130
rect 112 2106 146 2122
rect 112 114 146 130
rect 370 2106 404 2122
rect 370 114 404 130
rect -358 37 -342 71
rect -174 37 -158 71
rect -100 37 -84 71
rect 84 37 100 71
rect 158 37 174 71
rect 342 37 358 71
rect -358 -71 -342 -37
rect -174 -71 -158 -37
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect 158 -71 174 -37
rect 342 -71 358 -37
rect -404 -130 -370 -114
rect -404 -2122 -370 -2106
rect -146 -130 -112 -114
rect -146 -2122 -112 -2106
rect 112 -130 146 -114
rect 112 -2122 146 -2106
rect 370 -130 404 -114
rect 370 -2122 404 -2106
rect -358 -2199 -342 -2165
rect -174 -2199 -158 -2165
rect -100 -2199 -84 -2165
rect 84 -2199 100 -2165
rect 158 -2199 174 -2165
rect 342 -2199 358 -2165
rect -518 -2267 -484 -2205
rect 484 -2267 518 -2205
rect -518 -2301 -422 -2267
rect 422 -2301 518 -2267
<< viali >>
rect -342 2165 -174 2199
rect -84 2165 84 2199
rect 174 2165 342 2199
rect -404 130 -370 2106
rect -146 130 -112 2106
rect 112 130 146 2106
rect 370 130 404 2106
rect -342 37 -174 71
rect -84 37 84 71
rect 174 37 342 71
rect -342 -71 -174 -37
rect -84 -71 84 -37
rect 174 -71 342 -37
rect -404 -2106 -370 -130
rect -146 -2106 -112 -130
rect 112 -2106 146 -130
rect 370 -2106 404 -130
rect -342 -2199 -174 -2165
rect -84 -2199 84 -2165
rect 174 -2199 342 -2165
<< metal1 >>
rect -354 2199 -162 2205
rect -354 2165 -342 2199
rect -174 2165 -162 2199
rect -354 2159 -162 2165
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect 162 2199 354 2205
rect 162 2165 174 2199
rect 342 2165 354 2199
rect 162 2159 354 2165
rect -410 2106 -364 2118
rect -410 130 -404 2106
rect -370 130 -364 2106
rect -410 118 -364 130
rect -152 2106 -106 2118
rect -152 130 -146 2106
rect -112 130 -106 2106
rect -152 118 -106 130
rect 106 2106 152 2118
rect 106 130 112 2106
rect 146 130 152 2106
rect 106 118 152 130
rect 364 2106 410 2118
rect 364 130 370 2106
rect 404 130 410 2106
rect 364 118 410 130
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect -410 -130 -364 -118
rect -410 -2106 -404 -130
rect -370 -2106 -364 -130
rect -410 -2118 -364 -2106
rect -152 -130 -106 -118
rect -152 -2106 -146 -130
rect -112 -2106 -106 -130
rect -152 -2118 -106 -2106
rect 106 -130 152 -118
rect 106 -2106 112 -130
rect 146 -2106 152 -130
rect 106 -2118 152 -2106
rect 364 -130 410 -118
rect 364 -2106 370 -130
rect 404 -2106 410 -130
rect 364 -2118 410 -2106
rect -354 -2165 -162 -2159
rect -354 -2199 -342 -2165
rect -174 -2199 -162 -2165
rect -354 -2205 -162 -2199
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
rect 162 -2165 354 -2159
rect 162 -2199 174 -2165
rect 342 -2199 354 -2165
rect 162 -2205 354 -2199
<< properties >>
string FIXED_BBOX -501 -2284 501 2284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
