magic
tech sky130A
magscale 1 2
timestamp 1729267537
<< pwell >>
rect -1825 -2210 1825 2210
<< nmoslvt >>
rect -1629 -2000 -29 2000
rect 29 -2000 1629 2000
<< ndiff >>
rect -1687 1988 -1629 2000
rect -1687 -1988 -1675 1988
rect -1641 -1988 -1629 1988
rect -1687 -2000 -1629 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 1629 1988 1687 2000
rect 1629 -1988 1641 1988
rect 1675 -1988 1687 1988
rect 1629 -2000 1687 -1988
<< ndiffc >>
rect -1675 -1988 -1641 1988
rect -17 -1988 17 1988
rect 1641 -1988 1675 1988
<< psubdiff >>
rect -1789 2140 -1693 2174
rect 1693 2140 1789 2174
rect -1789 2078 -1755 2140
rect 1755 2078 1789 2140
rect -1789 -2140 -1755 -2078
rect 1755 -2140 1789 -2078
rect -1789 -2174 -1693 -2140
rect 1693 -2174 1789 -2140
<< psubdiffcont >>
rect -1693 2140 1693 2174
rect -1789 -2078 -1755 2078
rect 1755 -2078 1789 2078
rect -1693 -2174 1693 -2140
<< poly >>
rect -1629 2072 -29 2088
rect -1629 2038 -1613 2072
rect -45 2038 -29 2072
rect -1629 2000 -29 2038
rect 29 2072 1629 2088
rect 29 2038 45 2072
rect 1613 2038 1629 2072
rect 29 2000 1629 2038
rect -1629 -2038 -29 -2000
rect -1629 -2072 -1613 -2038
rect -45 -2072 -29 -2038
rect -1629 -2088 -29 -2072
rect 29 -2038 1629 -2000
rect 29 -2072 45 -2038
rect 1613 -2072 1629 -2038
rect 29 -2088 1629 -2072
<< polycont >>
rect -1613 2038 -45 2072
rect 45 2038 1613 2072
rect -1613 -2072 -45 -2038
rect 45 -2072 1613 -2038
<< locali >>
rect -1789 2140 -1693 2174
rect 1693 2140 1789 2174
rect -1789 2078 -1755 2140
rect 1755 2078 1789 2140
rect -1629 2038 -1613 2072
rect -45 2038 -29 2072
rect 29 2038 45 2072
rect 1613 2038 1629 2072
rect -1675 1988 -1641 2004
rect -1675 -2004 -1641 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 1641 1988 1675 2004
rect 1641 -2004 1675 -1988
rect -1629 -2072 -1613 -2038
rect -45 -2072 -29 -2038
rect 29 -2072 45 -2038
rect 1613 -2072 1629 -2038
rect -1789 -2140 -1755 -2078
rect 1755 -2140 1789 -2078
rect -1789 -2174 -1693 -2140
rect 1693 -2174 1789 -2140
<< viali >>
rect -1613 2038 -45 2072
rect 45 2038 1613 2072
rect -1675 -1988 -1641 1988
rect -17 -1988 17 1988
rect 1641 -1988 1675 1988
rect -1613 -2072 -45 -2038
rect 45 -2072 1613 -2038
<< metal1 >>
rect -1625 2072 -33 2078
rect -1625 2038 -1613 2072
rect -45 2038 -33 2072
rect -1625 2032 -33 2038
rect 33 2072 1625 2078
rect 33 2038 45 2072
rect 1613 2038 1625 2072
rect 33 2032 1625 2038
rect -1681 1988 -1635 2000
rect -1681 -1988 -1675 1988
rect -1641 -1988 -1635 1988
rect -1681 -2000 -1635 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 1635 1988 1681 2000
rect 1635 -1988 1641 1988
rect 1675 -1988 1681 1988
rect 1635 -2000 1681 -1988
rect -1625 -2038 -33 -2032
rect -1625 -2072 -1613 -2038
rect -45 -2072 -33 -2038
rect -1625 -2078 -33 -2072
rect 33 -2038 1625 -2032
rect 33 -2072 45 -2038
rect 1613 -2072 1625 -2038
rect 33 -2078 1625 -2072
<< properties >>
string FIXED_BBOX -1772 -2157 1772 2157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 20.0 l 8.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
