magic
tech sky130A
magscale 1 2
timestamp 1730410385
<< metal3 >>
rect -2886 1012 2886 1040
rect -2886 -1012 2802 1012
rect 2866 -1012 2886 1012
rect -2886 -1040 2886 -1012
<< via3 >>
rect 2802 -1012 2866 1012
<< mimcap >>
rect -2846 960 2554 1000
rect -2846 -960 -2806 960
rect 2514 -960 2554 960
rect -2846 -1000 2554 -960
<< mimcapcontact >>
rect -2806 -960 2514 960
<< metal4 >>
rect 2786 1012 2882 1028
rect -2807 960 2515 961
rect -2807 -960 -2806 960
rect 2514 -960 2515 960
rect -2807 -961 2515 -960
rect 2786 -1012 2802 1012
rect 2866 -1012 2882 1012
rect 2786 -1028 2882 -1012
<< properties >>
string FIXED_BBOX -2886 -1040 2594 1040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 27.0 l 10.0 val 554.06 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
