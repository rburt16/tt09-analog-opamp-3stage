magic
tech sky130A
magscale 1 2
timestamp 1721842171
<< pwell >>
rect -296 -7373 296 7373
<< nmos >>
rect -100 5563 100 7163
rect -100 3745 100 5345
rect -100 1927 100 3527
rect -100 109 100 1709
rect -100 -1709 100 -109
rect -100 -3527 100 -1927
rect -100 -5345 100 -3745
rect -100 -7163 100 -5563
<< ndiff >>
rect -158 7151 -100 7163
rect -158 5575 -146 7151
rect -112 5575 -100 7151
rect -158 5563 -100 5575
rect 100 7151 158 7163
rect 100 5575 112 7151
rect 146 5575 158 7151
rect 100 5563 158 5575
rect -158 5333 -100 5345
rect -158 3757 -146 5333
rect -112 3757 -100 5333
rect -158 3745 -100 3757
rect 100 5333 158 5345
rect 100 3757 112 5333
rect 146 3757 158 5333
rect 100 3745 158 3757
rect -158 3515 -100 3527
rect -158 1939 -146 3515
rect -112 1939 -100 3515
rect -158 1927 -100 1939
rect 100 3515 158 3527
rect 100 1939 112 3515
rect 146 1939 158 3515
rect 100 1927 158 1939
rect -158 1697 -100 1709
rect -158 121 -146 1697
rect -112 121 -100 1697
rect -158 109 -100 121
rect 100 1697 158 1709
rect 100 121 112 1697
rect 146 121 158 1697
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1697 -146 -121
rect -112 -1697 -100 -121
rect -158 -1709 -100 -1697
rect 100 -121 158 -109
rect 100 -1697 112 -121
rect 146 -1697 158 -121
rect 100 -1709 158 -1697
rect -158 -1939 -100 -1927
rect -158 -3515 -146 -1939
rect -112 -3515 -100 -1939
rect -158 -3527 -100 -3515
rect 100 -1939 158 -1927
rect 100 -3515 112 -1939
rect 146 -3515 158 -1939
rect 100 -3527 158 -3515
rect -158 -3757 -100 -3745
rect -158 -5333 -146 -3757
rect -112 -5333 -100 -3757
rect -158 -5345 -100 -5333
rect 100 -3757 158 -3745
rect 100 -5333 112 -3757
rect 146 -5333 158 -3757
rect 100 -5345 158 -5333
rect -158 -5575 -100 -5563
rect -158 -7151 -146 -5575
rect -112 -7151 -100 -5575
rect -158 -7163 -100 -7151
rect 100 -5575 158 -5563
rect 100 -7151 112 -5575
rect 146 -7151 158 -5575
rect 100 -7163 158 -7151
<< ndiffc >>
rect -146 5575 -112 7151
rect 112 5575 146 7151
rect -146 3757 -112 5333
rect 112 3757 146 5333
rect -146 1939 -112 3515
rect 112 1939 146 3515
rect -146 121 -112 1697
rect 112 121 146 1697
rect -146 -1697 -112 -121
rect 112 -1697 146 -121
rect -146 -3515 -112 -1939
rect 112 -3515 146 -1939
rect -146 -5333 -112 -3757
rect 112 -5333 146 -3757
rect -146 -7151 -112 -5575
rect 112 -7151 146 -5575
<< psubdiff >>
rect -260 7303 -164 7337
rect 164 7303 260 7337
rect -260 7241 -226 7303
rect 226 7241 260 7303
rect -260 -7303 -226 -7241
rect 226 -7303 260 -7241
rect -260 -7337 -164 -7303
rect 164 -7337 260 -7303
<< psubdiffcont >>
rect -164 7303 164 7337
rect -260 -7241 -226 7241
rect 226 -7241 260 7241
rect -164 -7337 164 -7303
<< poly >>
rect -100 7235 100 7251
rect -100 7201 -84 7235
rect 84 7201 100 7235
rect -100 7163 100 7201
rect -100 5525 100 5563
rect -100 5491 -84 5525
rect 84 5491 100 5525
rect -100 5475 100 5491
rect -100 5417 100 5433
rect -100 5383 -84 5417
rect 84 5383 100 5417
rect -100 5345 100 5383
rect -100 3707 100 3745
rect -100 3673 -84 3707
rect 84 3673 100 3707
rect -100 3657 100 3673
rect -100 3599 100 3615
rect -100 3565 -84 3599
rect 84 3565 100 3599
rect -100 3527 100 3565
rect -100 1889 100 1927
rect -100 1855 -84 1889
rect 84 1855 100 1889
rect -100 1839 100 1855
rect -100 1781 100 1797
rect -100 1747 -84 1781
rect 84 1747 100 1781
rect -100 1709 100 1747
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1747 100 -1709
rect -100 -1781 -84 -1747
rect 84 -1781 100 -1747
rect -100 -1797 100 -1781
rect -100 -1855 100 -1839
rect -100 -1889 -84 -1855
rect 84 -1889 100 -1855
rect -100 -1927 100 -1889
rect -100 -3565 100 -3527
rect -100 -3599 -84 -3565
rect 84 -3599 100 -3565
rect -100 -3615 100 -3599
rect -100 -3673 100 -3657
rect -100 -3707 -84 -3673
rect 84 -3707 100 -3673
rect -100 -3745 100 -3707
rect -100 -5383 100 -5345
rect -100 -5417 -84 -5383
rect 84 -5417 100 -5383
rect -100 -5433 100 -5417
rect -100 -5491 100 -5475
rect -100 -5525 -84 -5491
rect 84 -5525 100 -5491
rect -100 -5563 100 -5525
rect -100 -7201 100 -7163
rect -100 -7235 -84 -7201
rect 84 -7235 100 -7201
rect -100 -7251 100 -7235
<< polycont >>
rect -84 7201 84 7235
rect -84 5491 84 5525
rect -84 5383 84 5417
rect -84 3673 84 3707
rect -84 3565 84 3599
rect -84 1855 84 1889
rect -84 1747 84 1781
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1781 84 -1747
rect -84 -1889 84 -1855
rect -84 -3599 84 -3565
rect -84 -3707 84 -3673
rect -84 -5417 84 -5383
rect -84 -5525 84 -5491
rect -84 -7235 84 -7201
<< locali >>
rect -260 7303 -164 7337
rect 164 7303 260 7337
rect -260 7241 -226 7303
rect 226 7241 260 7303
rect -100 7201 -84 7235
rect 84 7201 100 7235
rect -146 7151 -112 7167
rect -146 5559 -112 5575
rect 112 7151 146 7167
rect 112 5559 146 5575
rect -100 5491 -84 5525
rect 84 5491 100 5525
rect -100 5383 -84 5417
rect 84 5383 100 5417
rect -146 5333 -112 5349
rect -146 3741 -112 3757
rect 112 5333 146 5349
rect 112 3741 146 3757
rect -100 3673 -84 3707
rect 84 3673 100 3707
rect -100 3565 -84 3599
rect 84 3565 100 3599
rect -146 3515 -112 3531
rect -146 1923 -112 1939
rect 112 3515 146 3531
rect 112 1923 146 1939
rect -100 1855 -84 1889
rect 84 1855 100 1889
rect -100 1747 -84 1781
rect 84 1747 100 1781
rect -146 1697 -112 1713
rect -146 105 -112 121
rect 112 1697 146 1713
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1713 -112 -1697
rect 112 -121 146 -105
rect 112 -1713 146 -1697
rect -100 -1781 -84 -1747
rect 84 -1781 100 -1747
rect -100 -1889 -84 -1855
rect 84 -1889 100 -1855
rect -146 -1939 -112 -1923
rect -146 -3531 -112 -3515
rect 112 -1939 146 -1923
rect 112 -3531 146 -3515
rect -100 -3599 -84 -3565
rect 84 -3599 100 -3565
rect -100 -3707 -84 -3673
rect 84 -3707 100 -3673
rect -146 -3757 -112 -3741
rect -146 -5349 -112 -5333
rect 112 -3757 146 -3741
rect 112 -5349 146 -5333
rect -100 -5417 -84 -5383
rect 84 -5417 100 -5383
rect -100 -5525 -84 -5491
rect 84 -5525 100 -5491
rect -146 -5575 -112 -5559
rect -146 -7167 -112 -7151
rect 112 -5575 146 -5559
rect 112 -7167 146 -7151
rect -100 -7235 -84 -7201
rect 84 -7235 100 -7201
rect -260 -7303 -226 -7241
rect 226 -7303 260 -7241
rect -260 -7337 -164 -7303
rect 164 -7337 260 -7303
<< viali >>
rect -84 7201 84 7235
rect -146 5575 -112 7151
rect 112 5575 146 7151
rect -84 5491 84 5525
rect -84 5383 84 5417
rect -146 3757 -112 5333
rect 112 3757 146 5333
rect -84 3673 84 3707
rect -84 3565 84 3599
rect -146 1939 -112 3515
rect 112 1939 146 3515
rect -84 1855 84 1889
rect -84 1747 84 1781
rect -146 121 -112 1697
rect 112 121 146 1697
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1697 -112 -121
rect 112 -1697 146 -121
rect -84 -1781 84 -1747
rect -84 -1889 84 -1855
rect -146 -3515 -112 -1939
rect 112 -3515 146 -1939
rect -84 -3599 84 -3565
rect -84 -3707 84 -3673
rect -146 -5333 -112 -3757
rect 112 -5333 146 -3757
rect -84 -5417 84 -5383
rect -84 -5525 84 -5491
rect -146 -7151 -112 -5575
rect 112 -7151 146 -5575
rect -84 -7235 84 -7201
<< metal1 >>
rect -96 7235 96 7241
rect -96 7201 -84 7235
rect 84 7201 96 7235
rect -96 7195 96 7201
rect -152 7151 -106 7163
rect -152 5575 -146 7151
rect -112 5575 -106 7151
rect -152 5563 -106 5575
rect 106 7151 152 7163
rect 106 5575 112 7151
rect 146 5575 152 7151
rect 106 5563 152 5575
rect -96 5525 96 5531
rect -96 5491 -84 5525
rect 84 5491 96 5525
rect -96 5485 96 5491
rect -96 5417 96 5423
rect -96 5383 -84 5417
rect 84 5383 96 5417
rect -96 5377 96 5383
rect -152 5333 -106 5345
rect -152 3757 -146 5333
rect -112 3757 -106 5333
rect -152 3745 -106 3757
rect 106 5333 152 5345
rect 106 3757 112 5333
rect 146 3757 152 5333
rect 106 3745 152 3757
rect -96 3707 96 3713
rect -96 3673 -84 3707
rect 84 3673 96 3707
rect -96 3667 96 3673
rect -96 3599 96 3605
rect -96 3565 -84 3599
rect 84 3565 96 3599
rect -96 3559 96 3565
rect -152 3515 -106 3527
rect -152 1939 -146 3515
rect -112 1939 -106 3515
rect -152 1927 -106 1939
rect 106 3515 152 3527
rect 106 1939 112 3515
rect 146 1939 152 3515
rect 106 1927 152 1939
rect -96 1889 96 1895
rect -96 1855 -84 1889
rect 84 1855 96 1889
rect -96 1849 96 1855
rect -96 1781 96 1787
rect -96 1747 -84 1781
rect 84 1747 96 1781
rect -96 1741 96 1747
rect -152 1697 -106 1709
rect -152 121 -146 1697
rect -112 121 -106 1697
rect -152 109 -106 121
rect 106 1697 152 1709
rect 106 121 112 1697
rect 146 121 152 1697
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -1697 -146 -121
rect -112 -1697 -106 -121
rect -152 -1709 -106 -1697
rect 106 -121 152 -109
rect 106 -1697 112 -121
rect 146 -1697 152 -121
rect 106 -1709 152 -1697
rect -96 -1747 96 -1741
rect -96 -1781 -84 -1747
rect 84 -1781 96 -1747
rect -96 -1787 96 -1781
rect -96 -1855 96 -1849
rect -96 -1889 -84 -1855
rect 84 -1889 96 -1855
rect -96 -1895 96 -1889
rect -152 -1939 -106 -1927
rect -152 -3515 -146 -1939
rect -112 -3515 -106 -1939
rect -152 -3527 -106 -3515
rect 106 -1939 152 -1927
rect 106 -3515 112 -1939
rect 146 -3515 152 -1939
rect 106 -3527 152 -3515
rect -96 -3565 96 -3559
rect -96 -3599 -84 -3565
rect 84 -3599 96 -3565
rect -96 -3605 96 -3599
rect -96 -3673 96 -3667
rect -96 -3707 -84 -3673
rect 84 -3707 96 -3673
rect -96 -3713 96 -3707
rect -152 -3757 -106 -3745
rect -152 -5333 -146 -3757
rect -112 -5333 -106 -3757
rect -152 -5345 -106 -5333
rect 106 -3757 152 -3745
rect 106 -5333 112 -3757
rect 146 -5333 152 -3757
rect 106 -5345 152 -5333
rect -96 -5383 96 -5377
rect -96 -5417 -84 -5383
rect 84 -5417 96 -5383
rect -96 -5423 96 -5417
rect -96 -5491 96 -5485
rect -96 -5525 -84 -5491
rect 84 -5525 96 -5491
rect -96 -5531 96 -5525
rect -152 -5575 -106 -5563
rect -152 -7151 -146 -5575
rect -112 -7151 -106 -5575
rect -152 -7163 -106 -7151
rect 106 -5575 152 -5563
rect 106 -7151 112 -5575
rect 146 -7151 152 -5575
rect 106 -7163 152 -7151
rect -96 -7201 96 -7195
rect -96 -7235 -84 -7201
rect 84 -7235 96 -7201
rect -96 -7241 96 -7235
<< properties >>
string FIXED_BBOX -243 -7320 243 7320
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8.0 l 1.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
