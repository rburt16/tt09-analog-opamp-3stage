magic
tech sky130A
magscale 1 2
timestamp 1730139296
<< pwell >>
rect -596 -4191 596 4191
<< nmoslvt >>
rect -400 3381 400 3981
rect -400 2563 400 3163
rect -400 1745 400 2345
rect -400 927 400 1527
rect -400 109 400 709
rect -400 -709 400 -109
rect -400 -1527 400 -927
rect -400 -2345 400 -1745
rect -400 -3163 400 -2563
rect -400 -3981 400 -3381
<< ndiff >>
rect -458 3825 -400 3981
rect -458 3537 -446 3825
rect -412 3537 -400 3825
rect -458 3381 -400 3537
rect 400 3825 458 3981
rect 400 3537 412 3825
rect 446 3537 458 3825
rect 400 3381 458 3537
rect -458 3007 -400 3163
rect -458 2719 -446 3007
rect -412 2719 -400 3007
rect -458 2563 -400 2719
rect 400 3007 458 3163
rect 400 2719 412 3007
rect 446 2719 458 3007
rect 400 2563 458 2719
rect -458 2189 -400 2345
rect -458 1901 -446 2189
rect -412 1901 -400 2189
rect -458 1745 -400 1901
rect 400 2189 458 2345
rect 400 1901 412 2189
rect 446 1901 458 2189
rect 400 1745 458 1901
rect -458 1371 -400 1527
rect -458 1083 -446 1371
rect -412 1083 -400 1371
rect -458 927 -400 1083
rect 400 1371 458 1527
rect 400 1083 412 1371
rect 446 1083 458 1371
rect 400 927 458 1083
rect -458 553 -400 709
rect -458 265 -446 553
rect -412 265 -400 553
rect -458 109 -400 265
rect 400 553 458 709
rect 400 265 412 553
rect 446 265 458 553
rect 400 109 458 265
rect -458 -265 -400 -109
rect -458 -553 -446 -265
rect -412 -553 -400 -265
rect -458 -709 -400 -553
rect 400 -265 458 -109
rect 400 -553 412 -265
rect 446 -553 458 -265
rect 400 -709 458 -553
rect -458 -1083 -400 -927
rect -458 -1371 -446 -1083
rect -412 -1371 -400 -1083
rect -458 -1527 -400 -1371
rect 400 -1083 458 -927
rect 400 -1371 412 -1083
rect 446 -1371 458 -1083
rect 400 -1527 458 -1371
rect -458 -1901 -400 -1745
rect -458 -2189 -446 -1901
rect -412 -2189 -400 -1901
rect -458 -2345 -400 -2189
rect 400 -1901 458 -1745
rect 400 -2189 412 -1901
rect 446 -2189 458 -1901
rect 400 -2345 458 -2189
rect -458 -2719 -400 -2563
rect -458 -3007 -446 -2719
rect -412 -3007 -400 -2719
rect -458 -3163 -400 -3007
rect 400 -2719 458 -2563
rect 400 -3007 412 -2719
rect 446 -3007 458 -2719
rect 400 -3163 458 -3007
rect -458 -3537 -400 -3381
rect -458 -3825 -446 -3537
rect -412 -3825 -400 -3537
rect -458 -3981 -400 -3825
rect 400 -3537 458 -3381
rect 400 -3825 412 -3537
rect 446 -3825 458 -3537
rect 400 -3981 458 -3825
<< ndiffc >>
rect -446 3537 -412 3825
rect 412 3537 446 3825
rect -446 2719 -412 3007
rect 412 2719 446 3007
rect -446 1901 -412 2189
rect 412 1901 446 2189
rect -446 1083 -412 1371
rect 412 1083 446 1371
rect -446 265 -412 553
rect 412 265 446 553
rect -446 -553 -412 -265
rect 412 -553 446 -265
rect -446 -1371 -412 -1083
rect 412 -1371 446 -1083
rect -446 -2189 -412 -1901
rect 412 -2189 446 -1901
rect -446 -3007 -412 -2719
rect 412 -3007 446 -2719
rect -446 -3825 -412 -3537
rect 412 -3825 446 -3537
<< psubdiff >>
rect -560 4121 -232 4155
rect 232 4121 560 4155
rect -560 2030 -526 4121
rect 526 2030 560 4121
rect -560 -4121 -526 -2030
rect 526 -4121 560 -2030
rect -560 -4155 -232 -4121
rect 232 -4155 560 -4121
<< psubdiffcont >>
rect -232 4121 232 4155
rect -560 -2030 -526 2030
rect 526 -2030 560 2030
rect -232 -4155 232 -4121
<< poly >>
rect -208 4053 208 4069
rect -208 4036 -192 4053
rect -400 4019 -192 4036
rect 192 4036 208 4053
rect 192 4019 400 4036
rect -400 3981 400 4019
rect -400 3343 400 3381
rect -400 3326 -192 3343
rect -208 3309 -192 3326
rect 192 3326 400 3343
rect 192 3309 208 3326
rect -208 3293 208 3309
rect -208 3235 208 3251
rect -208 3218 -192 3235
rect -400 3201 -192 3218
rect 192 3218 208 3235
rect 192 3201 400 3218
rect -400 3163 400 3201
rect -400 2525 400 2563
rect -400 2508 -192 2525
rect -208 2491 -192 2508
rect 192 2508 400 2525
rect 192 2491 208 2508
rect -208 2475 208 2491
rect -208 2417 208 2433
rect -208 2400 -192 2417
rect -400 2383 -192 2400
rect 192 2400 208 2417
rect 192 2383 400 2400
rect -400 2345 400 2383
rect -400 1707 400 1745
rect -400 1690 -192 1707
rect -208 1673 -192 1690
rect 192 1690 400 1707
rect 192 1673 208 1690
rect -208 1657 208 1673
rect -208 1599 208 1615
rect -208 1582 -192 1599
rect -400 1565 -192 1582
rect 192 1582 208 1599
rect 192 1565 400 1582
rect -400 1527 400 1565
rect -400 889 400 927
rect -400 872 -192 889
rect -208 855 -192 872
rect 192 872 400 889
rect 192 855 208 872
rect -208 839 208 855
rect -208 781 208 797
rect -208 764 -192 781
rect -400 747 -192 764
rect 192 764 208 781
rect 192 747 400 764
rect -400 709 400 747
rect -400 71 400 109
rect -400 54 -192 71
rect -208 37 -192 54
rect 192 54 400 71
rect 192 37 208 54
rect -208 21 208 37
rect -208 -37 208 -21
rect -208 -54 -192 -37
rect -400 -71 -192 -54
rect 192 -54 208 -37
rect 192 -71 400 -54
rect -400 -109 400 -71
rect -400 -747 400 -709
rect -400 -764 -192 -747
rect -208 -781 -192 -764
rect 192 -764 400 -747
rect 192 -781 208 -764
rect -208 -797 208 -781
rect -208 -855 208 -839
rect -208 -872 -192 -855
rect -400 -889 -192 -872
rect 192 -872 208 -855
rect 192 -889 400 -872
rect -400 -927 400 -889
rect -400 -1565 400 -1527
rect -400 -1582 -192 -1565
rect -208 -1599 -192 -1582
rect 192 -1582 400 -1565
rect 192 -1599 208 -1582
rect -208 -1615 208 -1599
rect -208 -1673 208 -1657
rect -208 -1690 -192 -1673
rect -400 -1707 -192 -1690
rect 192 -1690 208 -1673
rect 192 -1707 400 -1690
rect -400 -1745 400 -1707
rect -400 -2383 400 -2345
rect -400 -2400 -192 -2383
rect -208 -2417 -192 -2400
rect 192 -2400 400 -2383
rect 192 -2417 208 -2400
rect -208 -2433 208 -2417
rect -208 -2491 208 -2475
rect -208 -2508 -192 -2491
rect -400 -2525 -192 -2508
rect 192 -2508 208 -2491
rect 192 -2525 400 -2508
rect -400 -2563 400 -2525
rect -400 -3201 400 -3163
rect -400 -3218 -192 -3201
rect -208 -3235 -192 -3218
rect 192 -3218 400 -3201
rect 192 -3235 208 -3218
rect -208 -3251 208 -3235
rect -208 -3309 208 -3293
rect -208 -3326 -192 -3309
rect -400 -3343 -192 -3326
rect 192 -3326 208 -3309
rect 192 -3343 400 -3326
rect -400 -3381 400 -3343
rect -400 -4019 400 -3981
rect -400 -4036 -192 -4019
rect -208 -4053 -192 -4036
rect 192 -4036 400 -4019
rect 192 -4053 208 -4036
rect -208 -4069 208 -4053
<< polycont >>
rect -192 4019 192 4053
rect -192 3309 192 3343
rect -192 3201 192 3235
rect -192 2491 192 2525
rect -192 2383 192 2417
rect -192 1673 192 1707
rect -192 1565 192 1599
rect -192 855 192 889
rect -192 747 192 781
rect -192 37 192 71
rect -192 -71 192 -37
rect -192 -781 192 -747
rect -192 -889 192 -855
rect -192 -1599 192 -1565
rect -192 -1707 192 -1673
rect -192 -2417 192 -2383
rect -192 -2525 192 -2491
rect -192 -3235 192 -3201
rect -192 -3343 192 -3309
rect -192 -4053 192 -4019
<< locali >>
rect -560 4121 -263 4155
rect 263 4121 560 4155
rect -560 2061 -526 4121
rect -446 3825 -412 3841
rect -446 3521 -412 3537
rect 412 3825 446 3841
rect 412 3521 446 3537
rect -446 3007 -412 3023
rect -446 2703 -412 2719
rect 412 3007 446 3023
rect 412 2703 446 2719
rect -446 2189 -412 2205
rect -446 1885 -412 1901
rect 412 2189 446 2205
rect 412 1885 446 1901
rect 526 2061 560 4121
rect -446 1371 -412 1387
rect -446 1067 -412 1083
rect 412 1371 446 1387
rect 412 1067 446 1083
rect -446 553 -412 569
rect -446 249 -412 265
rect 412 553 446 569
rect 412 249 446 265
rect -446 -265 -412 -249
rect -446 -569 -412 -553
rect 412 -265 446 -249
rect 412 -569 446 -553
rect -446 -1083 -412 -1067
rect -446 -1387 -412 -1371
rect 412 -1083 446 -1067
rect 412 -1387 446 -1371
rect -560 -4121 -526 -2061
rect -446 -1901 -412 -1885
rect -446 -2205 -412 -2189
rect 412 -1901 446 -1885
rect 412 -2205 446 -2189
rect -446 -2719 -412 -2703
rect -446 -3023 -412 -3007
rect 412 -2719 446 -2703
rect 412 -3023 446 -3007
rect -446 -3537 -412 -3521
rect -446 -3841 -412 -3825
rect 412 -3537 446 -3521
rect 412 -3841 446 -3825
rect 526 -4121 560 -2061
rect -560 -4155 -263 -4121
rect 263 -4155 560 -4121
<< viali >>
rect -263 4121 -232 4155
rect -232 4121 232 4155
rect 232 4121 263 4155
rect -384 4019 -192 4053
rect -192 4019 192 4053
rect 192 4019 384 4053
rect -446 3537 -412 3825
rect 412 3537 446 3825
rect -384 3309 -192 3343
rect -192 3309 192 3343
rect 192 3309 384 3343
rect -384 3201 -192 3235
rect -192 3201 192 3235
rect 192 3201 384 3235
rect -446 2719 -412 3007
rect 412 2719 446 3007
rect -384 2491 -192 2525
rect -192 2491 192 2525
rect 192 2491 384 2525
rect -384 2383 -192 2417
rect -192 2383 192 2417
rect 192 2383 384 2417
rect -560 2030 -526 2061
rect -560 -2030 -526 2030
rect -446 1901 -412 2189
rect 412 1901 446 2189
rect 526 2030 560 2061
rect -384 1673 -192 1707
rect -192 1673 192 1707
rect 192 1673 384 1707
rect -384 1565 -192 1599
rect -192 1565 192 1599
rect 192 1565 384 1599
rect -446 1083 -412 1371
rect 412 1083 446 1371
rect -384 855 -192 889
rect -192 855 192 889
rect 192 855 384 889
rect -384 747 -192 781
rect -192 747 192 781
rect 192 747 384 781
rect -446 265 -412 553
rect 412 265 446 553
rect -384 37 -192 71
rect -192 37 192 71
rect 192 37 384 71
rect -384 -71 -192 -37
rect -192 -71 192 -37
rect 192 -71 384 -37
rect -446 -553 -412 -265
rect 412 -553 446 -265
rect -384 -781 -192 -747
rect -192 -781 192 -747
rect 192 -781 384 -747
rect -384 -889 -192 -855
rect -192 -889 192 -855
rect 192 -889 384 -855
rect -446 -1371 -412 -1083
rect 412 -1371 446 -1083
rect -384 -1599 -192 -1565
rect -192 -1599 192 -1565
rect 192 -1599 384 -1565
rect -384 -1707 -192 -1673
rect -192 -1707 192 -1673
rect 192 -1707 384 -1673
rect -560 -2061 -526 -2030
rect -446 -2189 -412 -1901
rect 412 -2189 446 -1901
rect 526 -2030 560 2030
rect 526 -2061 560 -2030
rect -384 -2417 -192 -2383
rect -192 -2417 192 -2383
rect 192 -2417 384 -2383
rect -384 -2525 -192 -2491
rect -192 -2525 192 -2491
rect 192 -2525 384 -2491
rect -446 -3007 -412 -2719
rect 412 -3007 446 -2719
rect -384 -3235 -192 -3201
rect -192 -3235 192 -3201
rect 192 -3235 384 -3201
rect -384 -3343 -192 -3309
rect -192 -3343 192 -3309
rect 192 -3343 384 -3309
rect -446 -3825 -412 -3537
rect 412 -3825 446 -3537
rect -384 -4053 -192 -4019
rect -192 -4053 192 -4019
rect 192 -4053 384 -4019
rect -263 -4155 -232 -4121
rect -232 -4155 232 -4121
rect 232 -4155 263 -4121
<< metal1 >>
rect -275 4155 275 4161
rect -275 4121 -263 4155
rect 263 4121 275 4155
rect -275 4115 275 4121
rect -396 4053 396 4059
rect -396 4019 -384 4053
rect 384 4019 396 4053
rect -396 4013 396 4019
rect -452 3825 -406 3837
rect -452 3537 -446 3825
rect -412 3537 -406 3825
rect -452 3525 -406 3537
rect 406 3825 452 3837
rect 406 3537 412 3825
rect 446 3537 452 3825
rect 406 3525 452 3537
rect -396 3343 396 3349
rect -396 3309 -384 3343
rect 384 3309 396 3343
rect -396 3303 396 3309
rect -396 3235 396 3241
rect -396 3201 -384 3235
rect 384 3201 396 3235
rect -396 3195 396 3201
rect -452 3007 -406 3019
rect -452 2719 -446 3007
rect -412 2719 -406 3007
rect -452 2707 -406 2719
rect 406 3007 452 3019
rect 406 2719 412 3007
rect 446 2719 452 3007
rect 406 2707 452 2719
rect -396 2525 396 2531
rect -396 2491 -384 2525
rect 384 2491 396 2525
rect -396 2485 396 2491
rect -396 2417 396 2423
rect -396 2383 -384 2417
rect 384 2383 396 2417
rect -396 2377 396 2383
rect -452 2189 -406 2201
rect -566 2061 -520 2073
rect -566 -2061 -560 2061
rect -526 -2061 -520 2061
rect -452 1901 -446 2189
rect -412 1901 -406 2189
rect -452 1889 -406 1901
rect 406 2189 452 2201
rect 406 1901 412 2189
rect 446 1901 452 2189
rect 406 1889 452 1901
rect 520 2061 566 2073
rect -396 1707 396 1713
rect -396 1673 -384 1707
rect 384 1673 396 1707
rect -396 1667 396 1673
rect -396 1599 396 1605
rect -396 1565 -384 1599
rect 384 1565 396 1599
rect -396 1559 396 1565
rect -452 1371 -406 1383
rect -452 1083 -446 1371
rect -412 1083 -406 1371
rect -452 1071 -406 1083
rect 406 1371 452 1383
rect 406 1083 412 1371
rect 446 1083 452 1371
rect 406 1071 452 1083
rect -396 889 396 895
rect -396 855 -384 889
rect 384 855 396 889
rect -396 849 396 855
rect -396 781 396 787
rect -396 747 -384 781
rect 384 747 396 781
rect -396 741 396 747
rect -452 553 -406 565
rect -452 265 -446 553
rect -412 265 -406 553
rect -452 253 -406 265
rect 406 553 452 565
rect 406 265 412 553
rect 446 265 452 553
rect 406 253 452 265
rect -396 71 396 77
rect -396 37 -384 71
rect 384 37 396 71
rect -396 31 396 37
rect -396 -37 396 -31
rect -396 -71 -384 -37
rect 384 -71 396 -37
rect -396 -77 396 -71
rect -452 -265 -406 -253
rect -452 -553 -446 -265
rect -412 -553 -406 -265
rect -452 -565 -406 -553
rect 406 -265 452 -253
rect 406 -553 412 -265
rect 446 -553 452 -265
rect 406 -565 452 -553
rect -396 -747 396 -741
rect -396 -781 -384 -747
rect 384 -781 396 -747
rect -396 -787 396 -781
rect -396 -855 396 -849
rect -396 -889 -384 -855
rect 384 -889 396 -855
rect -396 -895 396 -889
rect -452 -1083 -406 -1071
rect -452 -1371 -446 -1083
rect -412 -1371 -406 -1083
rect -452 -1383 -406 -1371
rect 406 -1083 452 -1071
rect 406 -1371 412 -1083
rect 446 -1371 452 -1083
rect 406 -1383 452 -1371
rect -396 -1565 396 -1559
rect -396 -1599 -384 -1565
rect 384 -1599 396 -1565
rect -396 -1605 396 -1599
rect -396 -1673 396 -1667
rect -396 -1707 -384 -1673
rect 384 -1707 396 -1673
rect -396 -1713 396 -1707
rect -566 -2073 -520 -2061
rect -452 -1901 -406 -1889
rect -452 -2189 -446 -1901
rect -412 -2189 -406 -1901
rect -452 -2201 -406 -2189
rect 406 -1901 452 -1889
rect 406 -2189 412 -1901
rect 446 -2189 452 -1901
rect 520 -2061 526 2061
rect 560 -2061 566 2061
rect 520 -2073 566 -2061
rect 406 -2201 452 -2189
rect -396 -2383 396 -2377
rect -396 -2417 -384 -2383
rect 384 -2417 396 -2383
rect -396 -2423 396 -2417
rect -396 -2491 396 -2485
rect -396 -2525 -384 -2491
rect 384 -2525 396 -2491
rect -396 -2531 396 -2525
rect -452 -2719 -406 -2707
rect -452 -3007 -446 -2719
rect -412 -3007 -406 -2719
rect -452 -3019 -406 -3007
rect 406 -2719 452 -2707
rect 406 -3007 412 -2719
rect 446 -3007 452 -2719
rect 406 -3019 452 -3007
rect -396 -3201 396 -3195
rect -396 -3235 -384 -3201
rect 384 -3235 396 -3201
rect -396 -3241 396 -3235
rect -396 -3309 396 -3303
rect -396 -3343 -384 -3309
rect 384 -3343 396 -3309
rect -396 -3349 396 -3343
rect -452 -3537 -406 -3525
rect -452 -3825 -446 -3537
rect -412 -3825 -406 -3537
rect -452 -3837 -406 -3825
rect 406 -3537 452 -3525
rect 406 -3825 412 -3537
rect 446 -3825 452 -3537
rect 406 -3837 452 -3825
rect -396 -4019 396 -4013
rect -396 -4053 -384 -4019
rect 384 -4053 396 -4019
rect -396 -4059 396 -4053
rect -275 -4121 275 -4115
rect -275 -4155 -263 -4121
rect 263 -4155 275 -4121
rect -275 -4161 275 -4155
<< properties >>
string FIXED_BBOX -543 -4138 543 4138
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3.0 l 4.0 m 10 nf 1 diffcov 50 polycov 50 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 50 rlcov 50 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 50 viadrn 50 viagate 100 viagb 50 viagr 50 viagl 50 viagt 50
<< end >>
