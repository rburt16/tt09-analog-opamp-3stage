magic
tech sky130A
magscale 1 2
timestamp 1727972425
<< nwell >>
rect -3335 -2219 3335 2219
<< pmoslvt >>
rect -3139 -2000 -2999 2000
rect -2941 -2000 -2801 2000
rect -2743 -2000 -2603 2000
rect -2545 -2000 -2405 2000
rect -2347 -2000 -2207 2000
rect -2149 -2000 -2009 2000
rect -1951 -2000 -1811 2000
rect -1753 -2000 -1613 2000
rect -1555 -2000 -1415 2000
rect -1357 -2000 -1217 2000
rect -1159 -2000 -1019 2000
rect -961 -2000 -821 2000
rect -763 -2000 -623 2000
rect -565 -2000 -425 2000
rect -367 -2000 -227 2000
rect -169 -2000 -29 2000
rect 29 -2000 169 2000
rect 227 -2000 367 2000
rect 425 -2000 565 2000
rect 623 -2000 763 2000
rect 821 -2000 961 2000
rect 1019 -2000 1159 2000
rect 1217 -2000 1357 2000
rect 1415 -2000 1555 2000
rect 1613 -2000 1753 2000
rect 1811 -2000 1951 2000
rect 2009 -2000 2149 2000
rect 2207 -2000 2347 2000
rect 2405 -2000 2545 2000
rect 2603 -2000 2743 2000
rect 2801 -2000 2941 2000
rect 2999 -2000 3139 2000
<< pdiff >>
rect -3197 1988 -3139 2000
rect -3197 -1988 -3185 1988
rect -3151 -1988 -3139 1988
rect -3197 -2000 -3139 -1988
rect -2999 1988 -2941 2000
rect -2999 -1988 -2987 1988
rect -2953 -1988 -2941 1988
rect -2999 -2000 -2941 -1988
rect -2801 1988 -2743 2000
rect -2801 -1988 -2789 1988
rect -2755 -1988 -2743 1988
rect -2801 -2000 -2743 -1988
rect -2603 1988 -2545 2000
rect -2603 -1988 -2591 1988
rect -2557 -1988 -2545 1988
rect -2603 -2000 -2545 -1988
rect -2405 1988 -2347 2000
rect -2405 -1988 -2393 1988
rect -2359 -1988 -2347 1988
rect -2405 -2000 -2347 -1988
rect -2207 1988 -2149 2000
rect -2207 -1988 -2195 1988
rect -2161 -1988 -2149 1988
rect -2207 -2000 -2149 -1988
rect -2009 1988 -1951 2000
rect -2009 -1988 -1997 1988
rect -1963 -1988 -1951 1988
rect -2009 -2000 -1951 -1988
rect -1811 1988 -1753 2000
rect -1811 -1988 -1799 1988
rect -1765 -1988 -1753 1988
rect -1811 -2000 -1753 -1988
rect -1613 1988 -1555 2000
rect -1613 -1988 -1601 1988
rect -1567 -1988 -1555 1988
rect -1613 -2000 -1555 -1988
rect -1415 1988 -1357 2000
rect -1415 -1988 -1403 1988
rect -1369 -1988 -1357 1988
rect -1415 -2000 -1357 -1988
rect -1217 1988 -1159 2000
rect -1217 -1988 -1205 1988
rect -1171 -1988 -1159 1988
rect -1217 -2000 -1159 -1988
rect -1019 1988 -961 2000
rect -1019 -1988 -1007 1988
rect -973 -1988 -961 1988
rect -1019 -2000 -961 -1988
rect -821 1988 -763 2000
rect -821 -1988 -809 1988
rect -775 -1988 -763 1988
rect -821 -2000 -763 -1988
rect -623 1988 -565 2000
rect -623 -1988 -611 1988
rect -577 -1988 -565 1988
rect -623 -2000 -565 -1988
rect -425 1988 -367 2000
rect -425 -1988 -413 1988
rect -379 -1988 -367 1988
rect -425 -2000 -367 -1988
rect -227 1988 -169 2000
rect -227 -1988 -215 1988
rect -181 -1988 -169 1988
rect -227 -2000 -169 -1988
rect -29 1988 29 2000
rect -29 -1988 -17 1988
rect 17 -1988 29 1988
rect -29 -2000 29 -1988
rect 169 1988 227 2000
rect 169 -1988 181 1988
rect 215 -1988 227 1988
rect 169 -2000 227 -1988
rect 367 1988 425 2000
rect 367 -1988 379 1988
rect 413 -1988 425 1988
rect 367 -2000 425 -1988
rect 565 1988 623 2000
rect 565 -1988 577 1988
rect 611 -1988 623 1988
rect 565 -2000 623 -1988
rect 763 1988 821 2000
rect 763 -1988 775 1988
rect 809 -1988 821 1988
rect 763 -2000 821 -1988
rect 961 1988 1019 2000
rect 961 -1988 973 1988
rect 1007 -1988 1019 1988
rect 961 -2000 1019 -1988
rect 1159 1988 1217 2000
rect 1159 -1988 1171 1988
rect 1205 -1988 1217 1988
rect 1159 -2000 1217 -1988
rect 1357 1988 1415 2000
rect 1357 -1988 1369 1988
rect 1403 -1988 1415 1988
rect 1357 -2000 1415 -1988
rect 1555 1988 1613 2000
rect 1555 -1988 1567 1988
rect 1601 -1988 1613 1988
rect 1555 -2000 1613 -1988
rect 1753 1988 1811 2000
rect 1753 -1988 1765 1988
rect 1799 -1988 1811 1988
rect 1753 -2000 1811 -1988
rect 1951 1988 2009 2000
rect 1951 -1988 1963 1988
rect 1997 -1988 2009 1988
rect 1951 -2000 2009 -1988
rect 2149 1988 2207 2000
rect 2149 -1988 2161 1988
rect 2195 -1988 2207 1988
rect 2149 -2000 2207 -1988
rect 2347 1988 2405 2000
rect 2347 -1988 2359 1988
rect 2393 -1988 2405 1988
rect 2347 -2000 2405 -1988
rect 2545 1988 2603 2000
rect 2545 -1988 2557 1988
rect 2591 -1988 2603 1988
rect 2545 -2000 2603 -1988
rect 2743 1988 2801 2000
rect 2743 -1988 2755 1988
rect 2789 -1988 2801 1988
rect 2743 -2000 2801 -1988
rect 2941 1988 2999 2000
rect 2941 -1988 2953 1988
rect 2987 -1988 2999 1988
rect 2941 -2000 2999 -1988
rect 3139 1988 3197 2000
rect 3139 -1988 3151 1988
rect 3185 -1988 3197 1988
rect 3139 -2000 3197 -1988
<< pdiffc >>
rect -3185 -1988 -3151 1988
rect -2987 -1988 -2953 1988
rect -2789 -1988 -2755 1988
rect -2591 -1988 -2557 1988
rect -2393 -1988 -2359 1988
rect -2195 -1988 -2161 1988
rect -1997 -1988 -1963 1988
rect -1799 -1988 -1765 1988
rect -1601 -1988 -1567 1988
rect -1403 -1988 -1369 1988
rect -1205 -1988 -1171 1988
rect -1007 -1988 -973 1988
rect -809 -1988 -775 1988
rect -611 -1988 -577 1988
rect -413 -1988 -379 1988
rect -215 -1988 -181 1988
rect -17 -1988 17 1988
rect 181 -1988 215 1988
rect 379 -1988 413 1988
rect 577 -1988 611 1988
rect 775 -1988 809 1988
rect 973 -1988 1007 1988
rect 1171 -1988 1205 1988
rect 1369 -1988 1403 1988
rect 1567 -1988 1601 1988
rect 1765 -1988 1799 1988
rect 1963 -1988 1997 1988
rect 2161 -1988 2195 1988
rect 2359 -1988 2393 1988
rect 2557 -1988 2591 1988
rect 2755 -1988 2789 1988
rect 2953 -1988 2987 1988
rect 3151 -1988 3185 1988
<< nsubdiff >>
rect -3299 2149 -3203 2183
rect 3203 2149 3299 2183
rect -3299 2087 -3265 2149
rect 3265 2087 3299 2149
rect -3299 -2149 -3265 -2087
rect 3265 -2149 3299 -2087
rect -3299 -2183 -3203 -2149
rect 3203 -2183 3299 -2149
<< nsubdiffcont >>
rect -3203 2149 3203 2183
rect -3299 -2087 -3265 2087
rect 3265 -2087 3299 2087
rect -3203 -2183 3203 -2149
<< poly >>
rect -3139 2081 -2999 2097
rect -3139 2047 -3123 2081
rect -3015 2047 -2999 2081
rect -3139 2000 -2999 2047
rect -2941 2081 -2801 2097
rect -2941 2047 -2925 2081
rect -2817 2047 -2801 2081
rect -2941 2000 -2801 2047
rect -2743 2081 -2603 2097
rect -2743 2047 -2727 2081
rect -2619 2047 -2603 2081
rect -2743 2000 -2603 2047
rect -2545 2081 -2405 2097
rect -2545 2047 -2529 2081
rect -2421 2047 -2405 2081
rect -2545 2000 -2405 2047
rect -2347 2081 -2207 2097
rect -2347 2047 -2331 2081
rect -2223 2047 -2207 2081
rect -2347 2000 -2207 2047
rect -2149 2081 -2009 2097
rect -2149 2047 -2133 2081
rect -2025 2047 -2009 2081
rect -2149 2000 -2009 2047
rect -1951 2081 -1811 2097
rect -1951 2047 -1935 2081
rect -1827 2047 -1811 2081
rect -1951 2000 -1811 2047
rect -1753 2081 -1613 2097
rect -1753 2047 -1737 2081
rect -1629 2047 -1613 2081
rect -1753 2000 -1613 2047
rect -1555 2081 -1415 2097
rect -1555 2047 -1539 2081
rect -1431 2047 -1415 2081
rect -1555 2000 -1415 2047
rect -1357 2081 -1217 2097
rect -1357 2047 -1341 2081
rect -1233 2047 -1217 2081
rect -1357 2000 -1217 2047
rect -1159 2081 -1019 2097
rect -1159 2047 -1143 2081
rect -1035 2047 -1019 2081
rect -1159 2000 -1019 2047
rect -961 2081 -821 2097
rect -961 2047 -945 2081
rect -837 2047 -821 2081
rect -961 2000 -821 2047
rect -763 2081 -623 2097
rect -763 2047 -747 2081
rect -639 2047 -623 2081
rect -763 2000 -623 2047
rect -565 2081 -425 2097
rect -565 2047 -549 2081
rect -441 2047 -425 2081
rect -565 2000 -425 2047
rect -367 2081 -227 2097
rect -367 2047 -351 2081
rect -243 2047 -227 2081
rect -367 2000 -227 2047
rect -169 2081 -29 2097
rect -169 2047 -153 2081
rect -45 2047 -29 2081
rect -169 2000 -29 2047
rect 29 2081 169 2097
rect 29 2047 45 2081
rect 153 2047 169 2081
rect 29 2000 169 2047
rect 227 2081 367 2097
rect 227 2047 243 2081
rect 351 2047 367 2081
rect 227 2000 367 2047
rect 425 2081 565 2097
rect 425 2047 441 2081
rect 549 2047 565 2081
rect 425 2000 565 2047
rect 623 2081 763 2097
rect 623 2047 639 2081
rect 747 2047 763 2081
rect 623 2000 763 2047
rect 821 2081 961 2097
rect 821 2047 837 2081
rect 945 2047 961 2081
rect 821 2000 961 2047
rect 1019 2081 1159 2097
rect 1019 2047 1035 2081
rect 1143 2047 1159 2081
rect 1019 2000 1159 2047
rect 1217 2081 1357 2097
rect 1217 2047 1233 2081
rect 1341 2047 1357 2081
rect 1217 2000 1357 2047
rect 1415 2081 1555 2097
rect 1415 2047 1431 2081
rect 1539 2047 1555 2081
rect 1415 2000 1555 2047
rect 1613 2081 1753 2097
rect 1613 2047 1629 2081
rect 1737 2047 1753 2081
rect 1613 2000 1753 2047
rect 1811 2081 1951 2097
rect 1811 2047 1827 2081
rect 1935 2047 1951 2081
rect 1811 2000 1951 2047
rect 2009 2081 2149 2097
rect 2009 2047 2025 2081
rect 2133 2047 2149 2081
rect 2009 2000 2149 2047
rect 2207 2081 2347 2097
rect 2207 2047 2223 2081
rect 2331 2047 2347 2081
rect 2207 2000 2347 2047
rect 2405 2081 2545 2097
rect 2405 2047 2421 2081
rect 2529 2047 2545 2081
rect 2405 2000 2545 2047
rect 2603 2081 2743 2097
rect 2603 2047 2619 2081
rect 2727 2047 2743 2081
rect 2603 2000 2743 2047
rect 2801 2081 2941 2097
rect 2801 2047 2817 2081
rect 2925 2047 2941 2081
rect 2801 2000 2941 2047
rect 2999 2081 3139 2097
rect 2999 2047 3015 2081
rect 3123 2047 3139 2081
rect 2999 2000 3139 2047
rect -3139 -2047 -2999 -2000
rect -3139 -2081 -3123 -2047
rect -3015 -2081 -2999 -2047
rect -3139 -2097 -2999 -2081
rect -2941 -2047 -2801 -2000
rect -2941 -2081 -2925 -2047
rect -2817 -2081 -2801 -2047
rect -2941 -2097 -2801 -2081
rect -2743 -2047 -2603 -2000
rect -2743 -2081 -2727 -2047
rect -2619 -2081 -2603 -2047
rect -2743 -2097 -2603 -2081
rect -2545 -2047 -2405 -2000
rect -2545 -2081 -2529 -2047
rect -2421 -2081 -2405 -2047
rect -2545 -2097 -2405 -2081
rect -2347 -2047 -2207 -2000
rect -2347 -2081 -2331 -2047
rect -2223 -2081 -2207 -2047
rect -2347 -2097 -2207 -2081
rect -2149 -2047 -2009 -2000
rect -2149 -2081 -2133 -2047
rect -2025 -2081 -2009 -2047
rect -2149 -2097 -2009 -2081
rect -1951 -2047 -1811 -2000
rect -1951 -2081 -1935 -2047
rect -1827 -2081 -1811 -2047
rect -1951 -2097 -1811 -2081
rect -1753 -2047 -1613 -2000
rect -1753 -2081 -1737 -2047
rect -1629 -2081 -1613 -2047
rect -1753 -2097 -1613 -2081
rect -1555 -2047 -1415 -2000
rect -1555 -2081 -1539 -2047
rect -1431 -2081 -1415 -2047
rect -1555 -2097 -1415 -2081
rect -1357 -2047 -1217 -2000
rect -1357 -2081 -1341 -2047
rect -1233 -2081 -1217 -2047
rect -1357 -2097 -1217 -2081
rect -1159 -2047 -1019 -2000
rect -1159 -2081 -1143 -2047
rect -1035 -2081 -1019 -2047
rect -1159 -2097 -1019 -2081
rect -961 -2047 -821 -2000
rect -961 -2081 -945 -2047
rect -837 -2081 -821 -2047
rect -961 -2097 -821 -2081
rect -763 -2047 -623 -2000
rect -763 -2081 -747 -2047
rect -639 -2081 -623 -2047
rect -763 -2097 -623 -2081
rect -565 -2047 -425 -2000
rect -565 -2081 -549 -2047
rect -441 -2081 -425 -2047
rect -565 -2097 -425 -2081
rect -367 -2047 -227 -2000
rect -367 -2081 -351 -2047
rect -243 -2081 -227 -2047
rect -367 -2097 -227 -2081
rect -169 -2047 -29 -2000
rect -169 -2081 -153 -2047
rect -45 -2081 -29 -2047
rect -169 -2097 -29 -2081
rect 29 -2047 169 -2000
rect 29 -2081 45 -2047
rect 153 -2081 169 -2047
rect 29 -2097 169 -2081
rect 227 -2047 367 -2000
rect 227 -2081 243 -2047
rect 351 -2081 367 -2047
rect 227 -2097 367 -2081
rect 425 -2047 565 -2000
rect 425 -2081 441 -2047
rect 549 -2081 565 -2047
rect 425 -2097 565 -2081
rect 623 -2047 763 -2000
rect 623 -2081 639 -2047
rect 747 -2081 763 -2047
rect 623 -2097 763 -2081
rect 821 -2047 961 -2000
rect 821 -2081 837 -2047
rect 945 -2081 961 -2047
rect 821 -2097 961 -2081
rect 1019 -2047 1159 -2000
rect 1019 -2081 1035 -2047
rect 1143 -2081 1159 -2047
rect 1019 -2097 1159 -2081
rect 1217 -2047 1357 -2000
rect 1217 -2081 1233 -2047
rect 1341 -2081 1357 -2047
rect 1217 -2097 1357 -2081
rect 1415 -2047 1555 -2000
rect 1415 -2081 1431 -2047
rect 1539 -2081 1555 -2047
rect 1415 -2097 1555 -2081
rect 1613 -2047 1753 -2000
rect 1613 -2081 1629 -2047
rect 1737 -2081 1753 -2047
rect 1613 -2097 1753 -2081
rect 1811 -2047 1951 -2000
rect 1811 -2081 1827 -2047
rect 1935 -2081 1951 -2047
rect 1811 -2097 1951 -2081
rect 2009 -2047 2149 -2000
rect 2009 -2081 2025 -2047
rect 2133 -2081 2149 -2047
rect 2009 -2097 2149 -2081
rect 2207 -2047 2347 -2000
rect 2207 -2081 2223 -2047
rect 2331 -2081 2347 -2047
rect 2207 -2097 2347 -2081
rect 2405 -2047 2545 -2000
rect 2405 -2081 2421 -2047
rect 2529 -2081 2545 -2047
rect 2405 -2097 2545 -2081
rect 2603 -2047 2743 -2000
rect 2603 -2081 2619 -2047
rect 2727 -2081 2743 -2047
rect 2603 -2097 2743 -2081
rect 2801 -2047 2941 -2000
rect 2801 -2081 2817 -2047
rect 2925 -2081 2941 -2047
rect 2801 -2097 2941 -2081
rect 2999 -2047 3139 -2000
rect 2999 -2081 3015 -2047
rect 3123 -2081 3139 -2047
rect 2999 -2097 3139 -2081
<< polycont >>
rect -3123 2047 -3015 2081
rect -2925 2047 -2817 2081
rect -2727 2047 -2619 2081
rect -2529 2047 -2421 2081
rect -2331 2047 -2223 2081
rect -2133 2047 -2025 2081
rect -1935 2047 -1827 2081
rect -1737 2047 -1629 2081
rect -1539 2047 -1431 2081
rect -1341 2047 -1233 2081
rect -1143 2047 -1035 2081
rect -945 2047 -837 2081
rect -747 2047 -639 2081
rect -549 2047 -441 2081
rect -351 2047 -243 2081
rect -153 2047 -45 2081
rect 45 2047 153 2081
rect 243 2047 351 2081
rect 441 2047 549 2081
rect 639 2047 747 2081
rect 837 2047 945 2081
rect 1035 2047 1143 2081
rect 1233 2047 1341 2081
rect 1431 2047 1539 2081
rect 1629 2047 1737 2081
rect 1827 2047 1935 2081
rect 2025 2047 2133 2081
rect 2223 2047 2331 2081
rect 2421 2047 2529 2081
rect 2619 2047 2727 2081
rect 2817 2047 2925 2081
rect 3015 2047 3123 2081
rect -3123 -2081 -3015 -2047
rect -2925 -2081 -2817 -2047
rect -2727 -2081 -2619 -2047
rect -2529 -2081 -2421 -2047
rect -2331 -2081 -2223 -2047
rect -2133 -2081 -2025 -2047
rect -1935 -2081 -1827 -2047
rect -1737 -2081 -1629 -2047
rect -1539 -2081 -1431 -2047
rect -1341 -2081 -1233 -2047
rect -1143 -2081 -1035 -2047
rect -945 -2081 -837 -2047
rect -747 -2081 -639 -2047
rect -549 -2081 -441 -2047
rect -351 -2081 -243 -2047
rect -153 -2081 -45 -2047
rect 45 -2081 153 -2047
rect 243 -2081 351 -2047
rect 441 -2081 549 -2047
rect 639 -2081 747 -2047
rect 837 -2081 945 -2047
rect 1035 -2081 1143 -2047
rect 1233 -2081 1341 -2047
rect 1431 -2081 1539 -2047
rect 1629 -2081 1737 -2047
rect 1827 -2081 1935 -2047
rect 2025 -2081 2133 -2047
rect 2223 -2081 2331 -2047
rect 2421 -2081 2529 -2047
rect 2619 -2081 2727 -2047
rect 2817 -2081 2925 -2047
rect 3015 -2081 3123 -2047
<< locali >>
rect -3299 2149 -3203 2183
rect 3203 2149 3299 2183
rect -3299 2087 -3265 2149
rect 3265 2087 3299 2149
rect -3139 2047 -3123 2081
rect -3015 2047 -2999 2081
rect -2941 2047 -2925 2081
rect -2817 2047 -2801 2081
rect -2743 2047 -2727 2081
rect -2619 2047 -2603 2081
rect -2545 2047 -2529 2081
rect -2421 2047 -2405 2081
rect -2347 2047 -2331 2081
rect -2223 2047 -2207 2081
rect -2149 2047 -2133 2081
rect -2025 2047 -2009 2081
rect -1951 2047 -1935 2081
rect -1827 2047 -1811 2081
rect -1753 2047 -1737 2081
rect -1629 2047 -1613 2081
rect -1555 2047 -1539 2081
rect -1431 2047 -1415 2081
rect -1357 2047 -1341 2081
rect -1233 2047 -1217 2081
rect -1159 2047 -1143 2081
rect -1035 2047 -1019 2081
rect -961 2047 -945 2081
rect -837 2047 -821 2081
rect -763 2047 -747 2081
rect -639 2047 -623 2081
rect -565 2047 -549 2081
rect -441 2047 -425 2081
rect -367 2047 -351 2081
rect -243 2047 -227 2081
rect -169 2047 -153 2081
rect -45 2047 -29 2081
rect 29 2047 45 2081
rect 153 2047 169 2081
rect 227 2047 243 2081
rect 351 2047 367 2081
rect 425 2047 441 2081
rect 549 2047 565 2081
rect 623 2047 639 2081
rect 747 2047 763 2081
rect 821 2047 837 2081
rect 945 2047 961 2081
rect 1019 2047 1035 2081
rect 1143 2047 1159 2081
rect 1217 2047 1233 2081
rect 1341 2047 1357 2081
rect 1415 2047 1431 2081
rect 1539 2047 1555 2081
rect 1613 2047 1629 2081
rect 1737 2047 1753 2081
rect 1811 2047 1827 2081
rect 1935 2047 1951 2081
rect 2009 2047 2025 2081
rect 2133 2047 2149 2081
rect 2207 2047 2223 2081
rect 2331 2047 2347 2081
rect 2405 2047 2421 2081
rect 2529 2047 2545 2081
rect 2603 2047 2619 2081
rect 2727 2047 2743 2081
rect 2801 2047 2817 2081
rect 2925 2047 2941 2081
rect 2999 2047 3015 2081
rect 3123 2047 3139 2081
rect -3185 1988 -3151 2004
rect -3185 -2004 -3151 -1988
rect -2987 1988 -2953 2004
rect -2987 -2004 -2953 -1988
rect -2789 1988 -2755 2004
rect -2789 -2004 -2755 -1988
rect -2591 1988 -2557 2004
rect -2591 -2004 -2557 -1988
rect -2393 1988 -2359 2004
rect -2393 -2004 -2359 -1988
rect -2195 1988 -2161 2004
rect -2195 -2004 -2161 -1988
rect -1997 1988 -1963 2004
rect -1997 -2004 -1963 -1988
rect -1799 1988 -1765 2004
rect -1799 -2004 -1765 -1988
rect -1601 1988 -1567 2004
rect -1601 -2004 -1567 -1988
rect -1403 1988 -1369 2004
rect -1403 -2004 -1369 -1988
rect -1205 1988 -1171 2004
rect -1205 -2004 -1171 -1988
rect -1007 1988 -973 2004
rect -1007 -2004 -973 -1988
rect -809 1988 -775 2004
rect -809 -2004 -775 -1988
rect -611 1988 -577 2004
rect -611 -2004 -577 -1988
rect -413 1988 -379 2004
rect -413 -2004 -379 -1988
rect -215 1988 -181 2004
rect -215 -2004 -181 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 181 1988 215 2004
rect 181 -2004 215 -1988
rect 379 1988 413 2004
rect 379 -2004 413 -1988
rect 577 1988 611 2004
rect 577 -2004 611 -1988
rect 775 1988 809 2004
rect 775 -2004 809 -1988
rect 973 1988 1007 2004
rect 973 -2004 1007 -1988
rect 1171 1988 1205 2004
rect 1171 -2004 1205 -1988
rect 1369 1988 1403 2004
rect 1369 -2004 1403 -1988
rect 1567 1988 1601 2004
rect 1567 -2004 1601 -1988
rect 1765 1988 1799 2004
rect 1765 -2004 1799 -1988
rect 1963 1988 1997 2004
rect 1963 -2004 1997 -1988
rect 2161 1988 2195 2004
rect 2161 -2004 2195 -1988
rect 2359 1988 2393 2004
rect 2359 -2004 2393 -1988
rect 2557 1988 2591 2004
rect 2557 -2004 2591 -1988
rect 2755 1988 2789 2004
rect 2755 -2004 2789 -1988
rect 2953 1988 2987 2004
rect 2953 -2004 2987 -1988
rect 3151 1988 3185 2004
rect 3151 -2004 3185 -1988
rect -3139 -2081 -3123 -2047
rect -3015 -2081 -2999 -2047
rect -2941 -2081 -2925 -2047
rect -2817 -2081 -2801 -2047
rect -2743 -2081 -2727 -2047
rect -2619 -2081 -2603 -2047
rect -2545 -2081 -2529 -2047
rect -2421 -2081 -2405 -2047
rect -2347 -2081 -2331 -2047
rect -2223 -2081 -2207 -2047
rect -2149 -2081 -2133 -2047
rect -2025 -2081 -2009 -2047
rect -1951 -2081 -1935 -2047
rect -1827 -2081 -1811 -2047
rect -1753 -2081 -1737 -2047
rect -1629 -2081 -1613 -2047
rect -1555 -2081 -1539 -2047
rect -1431 -2081 -1415 -2047
rect -1357 -2081 -1341 -2047
rect -1233 -2081 -1217 -2047
rect -1159 -2081 -1143 -2047
rect -1035 -2081 -1019 -2047
rect -961 -2081 -945 -2047
rect -837 -2081 -821 -2047
rect -763 -2081 -747 -2047
rect -639 -2081 -623 -2047
rect -565 -2081 -549 -2047
rect -441 -2081 -425 -2047
rect -367 -2081 -351 -2047
rect -243 -2081 -227 -2047
rect -169 -2081 -153 -2047
rect -45 -2081 -29 -2047
rect 29 -2081 45 -2047
rect 153 -2081 169 -2047
rect 227 -2081 243 -2047
rect 351 -2081 367 -2047
rect 425 -2081 441 -2047
rect 549 -2081 565 -2047
rect 623 -2081 639 -2047
rect 747 -2081 763 -2047
rect 821 -2081 837 -2047
rect 945 -2081 961 -2047
rect 1019 -2081 1035 -2047
rect 1143 -2081 1159 -2047
rect 1217 -2081 1233 -2047
rect 1341 -2081 1357 -2047
rect 1415 -2081 1431 -2047
rect 1539 -2081 1555 -2047
rect 1613 -2081 1629 -2047
rect 1737 -2081 1753 -2047
rect 1811 -2081 1827 -2047
rect 1935 -2081 1951 -2047
rect 2009 -2081 2025 -2047
rect 2133 -2081 2149 -2047
rect 2207 -2081 2223 -2047
rect 2331 -2081 2347 -2047
rect 2405 -2081 2421 -2047
rect 2529 -2081 2545 -2047
rect 2603 -2081 2619 -2047
rect 2727 -2081 2743 -2047
rect 2801 -2081 2817 -2047
rect 2925 -2081 2941 -2047
rect 2999 -2081 3015 -2047
rect 3123 -2081 3139 -2047
rect -3299 -2149 -3265 -2087
rect 3265 -2149 3299 -2087
rect -3299 -2183 -3203 -2149
rect 3203 -2183 3299 -2149
<< viali >>
rect -3123 2047 -3015 2081
rect -2925 2047 -2817 2081
rect -2727 2047 -2619 2081
rect -2529 2047 -2421 2081
rect -2331 2047 -2223 2081
rect -2133 2047 -2025 2081
rect -1935 2047 -1827 2081
rect -1737 2047 -1629 2081
rect -1539 2047 -1431 2081
rect -1341 2047 -1233 2081
rect -1143 2047 -1035 2081
rect -945 2047 -837 2081
rect -747 2047 -639 2081
rect -549 2047 -441 2081
rect -351 2047 -243 2081
rect -153 2047 -45 2081
rect 45 2047 153 2081
rect 243 2047 351 2081
rect 441 2047 549 2081
rect 639 2047 747 2081
rect 837 2047 945 2081
rect 1035 2047 1143 2081
rect 1233 2047 1341 2081
rect 1431 2047 1539 2081
rect 1629 2047 1737 2081
rect 1827 2047 1935 2081
rect 2025 2047 2133 2081
rect 2223 2047 2331 2081
rect 2421 2047 2529 2081
rect 2619 2047 2727 2081
rect 2817 2047 2925 2081
rect 3015 2047 3123 2081
rect -3185 -1988 -3151 1988
rect -2987 -1988 -2953 1988
rect -2789 -1988 -2755 1988
rect -2591 -1988 -2557 1988
rect -2393 -1988 -2359 1988
rect -2195 -1988 -2161 1988
rect -1997 -1988 -1963 1988
rect -1799 -1988 -1765 1988
rect -1601 -1988 -1567 1988
rect -1403 -1988 -1369 1988
rect -1205 -1988 -1171 1988
rect -1007 -1988 -973 1988
rect -809 -1988 -775 1988
rect -611 -1988 -577 1988
rect -413 -1988 -379 1988
rect -215 -1988 -181 1988
rect -17 -1988 17 1988
rect 181 -1988 215 1988
rect 379 -1988 413 1988
rect 577 -1988 611 1988
rect 775 -1988 809 1988
rect 973 -1988 1007 1988
rect 1171 -1988 1205 1988
rect 1369 -1988 1403 1988
rect 1567 -1988 1601 1988
rect 1765 -1988 1799 1988
rect 1963 -1988 1997 1988
rect 2161 -1988 2195 1988
rect 2359 -1988 2393 1988
rect 2557 -1988 2591 1988
rect 2755 -1988 2789 1988
rect 2953 -1988 2987 1988
rect 3151 -1988 3185 1988
rect -3123 -2081 -3015 -2047
rect -2925 -2081 -2817 -2047
rect -2727 -2081 -2619 -2047
rect -2529 -2081 -2421 -2047
rect -2331 -2081 -2223 -2047
rect -2133 -2081 -2025 -2047
rect -1935 -2081 -1827 -2047
rect -1737 -2081 -1629 -2047
rect -1539 -2081 -1431 -2047
rect -1341 -2081 -1233 -2047
rect -1143 -2081 -1035 -2047
rect -945 -2081 -837 -2047
rect -747 -2081 -639 -2047
rect -549 -2081 -441 -2047
rect -351 -2081 -243 -2047
rect -153 -2081 -45 -2047
rect 45 -2081 153 -2047
rect 243 -2081 351 -2047
rect 441 -2081 549 -2047
rect 639 -2081 747 -2047
rect 837 -2081 945 -2047
rect 1035 -2081 1143 -2047
rect 1233 -2081 1341 -2047
rect 1431 -2081 1539 -2047
rect 1629 -2081 1737 -2047
rect 1827 -2081 1935 -2047
rect 2025 -2081 2133 -2047
rect 2223 -2081 2331 -2047
rect 2421 -2081 2529 -2047
rect 2619 -2081 2727 -2047
rect 2817 -2081 2925 -2047
rect 3015 -2081 3123 -2047
<< metal1 >>
rect -3135 2081 -3003 2087
rect -3135 2047 -3123 2081
rect -3015 2047 -3003 2081
rect -3135 2041 -3003 2047
rect -2937 2081 -2805 2087
rect -2937 2047 -2925 2081
rect -2817 2047 -2805 2081
rect -2937 2041 -2805 2047
rect -2739 2081 -2607 2087
rect -2739 2047 -2727 2081
rect -2619 2047 -2607 2081
rect -2739 2041 -2607 2047
rect -2541 2081 -2409 2087
rect -2541 2047 -2529 2081
rect -2421 2047 -2409 2081
rect -2541 2041 -2409 2047
rect -2343 2081 -2211 2087
rect -2343 2047 -2331 2081
rect -2223 2047 -2211 2081
rect -2343 2041 -2211 2047
rect -2145 2081 -2013 2087
rect -2145 2047 -2133 2081
rect -2025 2047 -2013 2081
rect -2145 2041 -2013 2047
rect -1947 2081 -1815 2087
rect -1947 2047 -1935 2081
rect -1827 2047 -1815 2081
rect -1947 2041 -1815 2047
rect -1749 2081 -1617 2087
rect -1749 2047 -1737 2081
rect -1629 2047 -1617 2081
rect -1749 2041 -1617 2047
rect -1551 2081 -1419 2087
rect -1551 2047 -1539 2081
rect -1431 2047 -1419 2081
rect -1551 2041 -1419 2047
rect -1353 2081 -1221 2087
rect -1353 2047 -1341 2081
rect -1233 2047 -1221 2081
rect -1353 2041 -1221 2047
rect -1155 2081 -1023 2087
rect -1155 2047 -1143 2081
rect -1035 2047 -1023 2081
rect -1155 2041 -1023 2047
rect -957 2081 -825 2087
rect -957 2047 -945 2081
rect -837 2047 -825 2081
rect -957 2041 -825 2047
rect -759 2081 -627 2087
rect -759 2047 -747 2081
rect -639 2047 -627 2081
rect -759 2041 -627 2047
rect -561 2081 -429 2087
rect -561 2047 -549 2081
rect -441 2047 -429 2081
rect -561 2041 -429 2047
rect -363 2081 -231 2087
rect -363 2047 -351 2081
rect -243 2047 -231 2081
rect -363 2041 -231 2047
rect -165 2081 -33 2087
rect -165 2047 -153 2081
rect -45 2047 -33 2081
rect -165 2041 -33 2047
rect 33 2081 165 2087
rect 33 2047 45 2081
rect 153 2047 165 2081
rect 33 2041 165 2047
rect 231 2081 363 2087
rect 231 2047 243 2081
rect 351 2047 363 2081
rect 231 2041 363 2047
rect 429 2081 561 2087
rect 429 2047 441 2081
rect 549 2047 561 2081
rect 429 2041 561 2047
rect 627 2081 759 2087
rect 627 2047 639 2081
rect 747 2047 759 2081
rect 627 2041 759 2047
rect 825 2081 957 2087
rect 825 2047 837 2081
rect 945 2047 957 2081
rect 825 2041 957 2047
rect 1023 2081 1155 2087
rect 1023 2047 1035 2081
rect 1143 2047 1155 2081
rect 1023 2041 1155 2047
rect 1221 2081 1353 2087
rect 1221 2047 1233 2081
rect 1341 2047 1353 2081
rect 1221 2041 1353 2047
rect 1419 2081 1551 2087
rect 1419 2047 1431 2081
rect 1539 2047 1551 2081
rect 1419 2041 1551 2047
rect 1617 2081 1749 2087
rect 1617 2047 1629 2081
rect 1737 2047 1749 2081
rect 1617 2041 1749 2047
rect 1815 2081 1947 2087
rect 1815 2047 1827 2081
rect 1935 2047 1947 2081
rect 1815 2041 1947 2047
rect 2013 2081 2145 2087
rect 2013 2047 2025 2081
rect 2133 2047 2145 2081
rect 2013 2041 2145 2047
rect 2211 2081 2343 2087
rect 2211 2047 2223 2081
rect 2331 2047 2343 2081
rect 2211 2041 2343 2047
rect 2409 2081 2541 2087
rect 2409 2047 2421 2081
rect 2529 2047 2541 2081
rect 2409 2041 2541 2047
rect 2607 2081 2739 2087
rect 2607 2047 2619 2081
rect 2727 2047 2739 2081
rect 2607 2041 2739 2047
rect 2805 2081 2937 2087
rect 2805 2047 2817 2081
rect 2925 2047 2937 2081
rect 2805 2041 2937 2047
rect 3003 2081 3135 2087
rect 3003 2047 3015 2081
rect 3123 2047 3135 2081
rect 3003 2041 3135 2047
rect -3191 1988 -3145 2000
rect -3191 -1988 -3185 1988
rect -3151 -1988 -3145 1988
rect -3191 -2000 -3145 -1988
rect -2993 1988 -2947 2000
rect -2993 -1988 -2987 1988
rect -2953 -1988 -2947 1988
rect -2993 -2000 -2947 -1988
rect -2795 1988 -2749 2000
rect -2795 -1988 -2789 1988
rect -2755 -1988 -2749 1988
rect -2795 -2000 -2749 -1988
rect -2597 1988 -2551 2000
rect -2597 -1988 -2591 1988
rect -2557 -1988 -2551 1988
rect -2597 -2000 -2551 -1988
rect -2399 1988 -2353 2000
rect -2399 -1988 -2393 1988
rect -2359 -1988 -2353 1988
rect -2399 -2000 -2353 -1988
rect -2201 1988 -2155 2000
rect -2201 -1988 -2195 1988
rect -2161 -1988 -2155 1988
rect -2201 -2000 -2155 -1988
rect -2003 1988 -1957 2000
rect -2003 -1988 -1997 1988
rect -1963 -1988 -1957 1988
rect -2003 -2000 -1957 -1988
rect -1805 1988 -1759 2000
rect -1805 -1988 -1799 1988
rect -1765 -1988 -1759 1988
rect -1805 -2000 -1759 -1988
rect -1607 1988 -1561 2000
rect -1607 -1988 -1601 1988
rect -1567 -1988 -1561 1988
rect -1607 -2000 -1561 -1988
rect -1409 1988 -1363 2000
rect -1409 -1988 -1403 1988
rect -1369 -1988 -1363 1988
rect -1409 -2000 -1363 -1988
rect -1211 1988 -1165 2000
rect -1211 -1988 -1205 1988
rect -1171 -1988 -1165 1988
rect -1211 -2000 -1165 -1988
rect -1013 1988 -967 2000
rect -1013 -1988 -1007 1988
rect -973 -1988 -967 1988
rect -1013 -2000 -967 -1988
rect -815 1988 -769 2000
rect -815 -1988 -809 1988
rect -775 -1988 -769 1988
rect -815 -2000 -769 -1988
rect -617 1988 -571 2000
rect -617 -1988 -611 1988
rect -577 -1988 -571 1988
rect -617 -2000 -571 -1988
rect -419 1988 -373 2000
rect -419 -1988 -413 1988
rect -379 -1988 -373 1988
rect -419 -2000 -373 -1988
rect -221 1988 -175 2000
rect -221 -1988 -215 1988
rect -181 -1988 -175 1988
rect -221 -2000 -175 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 175 1988 221 2000
rect 175 -1988 181 1988
rect 215 -1988 221 1988
rect 175 -2000 221 -1988
rect 373 1988 419 2000
rect 373 -1988 379 1988
rect 413 -1988 419 1988
rect 373 -2000 419 -1988
rect 571 1988 617 2000
rect 571 -1988 577 1988
rect 611 -1988 617 1988
rect 571 -2000 617 -1988
rect 769 1988 815 2000
rect 769 -1988 775 1988
rect 809 -1988 815 1988
rect 769 -2000 815 -1988
rect 967 1988 1013 2000
rect 967 -1988 973 1988
rect 1007 -1988 1013 1988
rect 967 -2000 1013 -1988
rect 1165 1988 1211 2000
rect 1165 -1988 1171 1988
rect 1205 -1988 1211 1988
rect 1165 -2000 1211 -1988
rect 1363 1988 1409 2000
rect 1363 -1988 1369 1988
rect 1403 -1988 1409 1988
rect 1363 -2000 1409 -1988
rect 1561 1988 1607 2000
rect 1561 -1988 1567 1988
rect 1601 -1988 1607 1988
rect 1561 -2000 1607 -1988
rect 1759 1988 1805 2000
rect 1759 -1988 1765 1988
rect 1799 -1988 1805 1988
rect 1759 -2000 1805 -1988
rect 1957 1988 2003 2000
rect 1957 -1988 1963 1988
rect 1997 -1988 2003 1988
rect 1957 -2000 2003 -1988
rect 2155 1988 2201 2000
rect 2155 -1988 2161 1988
rect 2195 -1988 2201 1988
rect 2155 -2000 2201 -1988
rect 2353 1988 2399 2000
rect 2353 -1988 2359 1988
rect 2393 -1988 2399 1988
rect 2353 -2000 2399 -1988
rect 2551 1988 2597 2000
rect 2551 -1988 2557 1988
rect 2591 -1988 2597 1988
rect 2551 -2000 2597 -1988
rect 2749 1988 2795 2000
rect 2749 -1988 2755 1988
rect 2789 -1988 2795 1988
rect 2749 -2000 2795 -1988
rect 2947 1988 2993 2000
rect 2947 -1988 2953 1988
rect 2987 -1988 2993 1988
rect 2947 -2000 2993 -1988
rect 3145 1988 3191 2000
rect 3145 -1988 3151 1988
rect 3185 -1988 3191 1988
rect 3145 -2000 3191 -1988
rect -3135 -2047 -3003 -2041
rect -3135 -2081 -3123 -2047
rect -3015 -2081 -3003 -2047
rect -3135 -2087 -3003 -2081
rect -2937 -2047 -2805 -2041
rect -2937 -2081 -2925 -2047
rect -2817 -2081 -2805 -2047
rect -2937 -2087 -2805 -2081
rect -2739 -2047 -2607 -2041
rect -2739 -2081 -2727 -2047
rect -2619 -2081 -2607 -2047
rect -2739 -2087 -2607 -2081
rect -2541 -2047 -2409 -2041
rect -2541 -2081 -2529 -2047
rect -2421 -2081 -2409 -2047
rect -2541 -2087 -2409 -2081
rect -2343 -2047 -2211 -2041
rect -2343 -2081 -2331 -2047
rect -2223 -2081 -2211 -2047
rect -2343 -2087 -2211 -2081
rect -2145 -2047 -2013 -2041
rect -2145 -2081 -2133 -2047
rect -2025 -2081 -2013 -2047
rect -2145 -2087 -2013 -2081
rect -1947 -2047 -1815 -2041
rect -1947 -2081 -1935 -2047
rect -1827 -2081 -1815 -2047
rect -1947 -2087 -1815 -2081
rect -1749 -2047 -1617 -2041
rect -1749 -2081 -1737 -2047
rect -1629 -2081 -1617 -2047
rect -1749 -2087 -1617 -2081
rect -1551 -2047 -1419 -2041
rect -1551 -2081 -1539 -2047
rect -1431 -2081 -1419 -2047
rect -1551 -2087 -1419 -2081
rect -1353 -2047 -1221 -2041
rect -1353 -2081 -1341 -2047
rect -1233 -2081 -1221 -2047
rect -1353 -2087 -1221 -2081
rect -1155 -2047 -1023 -2041
rect -1155 -2081 -1143 -2047
rect -1035 -2081 -1023 -2047
rect -1155 -2087 -1023 -2081
rect -957 -2047 -825 -2041
rect -957 -2081 -945 -2047
rect -837 -2081 -825 -2047
rect -957 -2087 -825 -2081
rect -759 -2047 -627 -2041
rect -759 -2081 -747 -2047
rect -639 -2081 -627 -2047
rect -759 -2087 -627 -2081
rect -561 -2047 -429 -2041
rect -561 -2081 -549 -2047
rect -441 -2081 -429 -2047
rect -561 -2087 -429 -2081
rect -363 -2047 -231 -2041
rect -363 -2081 -351 -2047
rect -243 -2081 -231 -2047
rect -363 -2087 -231 -2081
rect -165 -2047 -33 -2041
rect -165 -2081 -153 -2047
rect -45 -2081 -33 -2047
rect -165 -2087 -33 -2081
rect 33 -2047 165 -2041
rect 33 -2081 45 -2047
rect 153 -2081 165 -2047
rect 33 -2087 165 -2081
rect 231 -2047 363 -2041
rect 231 -2081 243 -2047
rect 351 -2081 363 -2047
rect 231 -2087 363 -2081
rect 429 -2047 561 -2041
rect 429 -2081 441 -2047
rect 549 -2081 561 -2047
rect 429 -2087 561 -2081
rect 627 -2047 759 -2041
rect 627 -2081 639 -2047
rect 747 -2081 759 -2047
rect 627 -2087 759 -2081
rect 825 -2047 957 -2041
rect 825 -2081 837 -2047
rect 945 -2081 957 -2047
rect 825 -2087 957 -2081
rect 1023 -2047 1155 -2041
rect 1023 -2081 1035 -2047
rect 1143 -2081 1155 -2047
rect 1023 -2087 1155 -2081
rect 1221 -2047 1353 -2041
rect 1221 -2081 1233 -2047
rect 1341 -2081 1353 -2047
rect 1221 -2087 1353 -2081
rect 1419 -2047 1551 -2041
rect 1419 -2081 1431 -2047
rect 1539 -2081 1551 -2047
rect 1419 -2087 1551 -2081
rect 1617 -2047 1749 -2041
rect 1617 -2081 1629 -2047
rect 1737 -2081 1749 -2047
rect 1617 -2087 1749 -2081
rect 1815 -2047 1947 -2041
rect 1815 -2081 1827 -2047
rect 1935 -2081 1947 -2047
rect 1815 -2087 1947 -2081
rect 2013 -2047 2145 -2041
rect 2013 -2081 2025 -2047
rect 2133 -2081 2145 -2047
rect 2013 -2087 2145 -2081
rect 2211 -2047 2343 -2041
rect 2211 -2081 2223 -2047
rect 2331 -2081 2343 -2047
rect 2211 -2087 2343 -2081
rect 2409 -2047 2541 -2041
rect 2409 -2081 2421 -2047
rect 2529 -2081 2541 -2047
rect 2409 -2087 2541 -2081
rect 2607 -2047 2739 -2041
rect 2607 -2081 2619 -2047
rect 2727 -2081 2739 -2047
rect 2607 -2087 2739 -2081
rect 2805 -2047 2937 -2041
rect 2805 -2081 2817 -2047
rect 2925 -2081 2937 -2047
rect 2805 -2087 2937 -2081
rect 3003 -2047 3135 -2041
rect 3003 -2081 3015 -2047
rect 3123 -2081 3135 -2047
rect 3003 -2087 3135 -2081
<< properties >>
string FIXED_BBOX -3282 -2166 3282 2166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 20.0 l 0.7 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
