magic
tech sky130A
magscale 1 2
timestamp 1728061155
<< metal3 >>
rect -13104 2812 -6732 2840
rect -13104 -2812 -6816 2812
rect -6752 -2812 -6732 2812
rect -13104 -2840 -6732 -2812
rect -6492 2812 -120 2840
rect -6492 -2812 -204 2812
rect -140 -2812 -120 2812
rect -6492 -2840 -120 -2812
rect 120 2812 6492 2840
rect 120 -2812 6408 2812
rect 6472 -2812 6492 2812
rect 120 -2840 6492 -2812
rect 6732 2812 13104 2840
rect 6732 -2812 13020 2812
rect 13084 -2812 13104 2812
rect 6732 -2840 13104 -2812
<< via3 >>
rect -6816 -2812 -6752 2812
rect -204 -2812 -140 2812
rect 6408 -2812 6472 2812
rect 13020 -2812 13084 2812
<< mimcap >>
rect -13064 2760 -7064 2800
rect -13064 -2760 -13024 2760
rect -7104 -2760 -7064 2760
rect -13064 -2800 -7064 -2760
rect -6452 2760 -452 2800
rect -6452 -2760 -6412 2760
rect -492 -2760 -452 2760
rect -6452 -2800 -452 -2760
rect 160 2760 6160 2800
rect 160 -2760 200 2760
rect 6120 -2760 6160 2760
rect 160 -2800 6160 -2760
rect 6772 2760 12772 2800
rect 6772 -2760 6812 2760
rect 12732 -2760 12772 2760
rect 6772 -2800 12772 -2760
<< mimcapcontact >>
rect -13024 -2760 -7104 2760
rect -6412 -2760 -492 2760
rect 200 -2760 6120 2760
rect 6812 -2760 12732 2760
<< metal4 >>
rect -6832 2812 -6736 2828
rect -13025 2760 -7103 2761
rect -13025 -2760 -13024 2760
rect -7104 -2760 -7103 2760
rect -13025 -2761 -7103 -2760
rect -6832 -2812 -6816 2812
rect -6752 -2812 -6736 2812
rect -220 2812 -124 2828
rect -6413 2760 -491 2761
rect -6413 -2760 -6412 2760
rect -492 -2760 -491 2760
rect -6413 -2761 -491 -2760
rect -6832 -2828 -6736 -2812
rect -220 -2812 -204 2812
rect -140 -2812 -124 2812
rect 6392 2812 6488 2828
rect 199 2760 6121 2761
rect 199 -2760 200 2760
rect 6120 -2760 6121 2760
rect 199 -2761 6121 -2760
rect -220 -2828 -124 -2812
rect 6392 -2812 6408 2812
rect 6472 -2812 6488 2812
rect 13004 2812 13100 2828
rect 6811 2760 12733 2761
rect 6811 -2760 6812 2760
rect 12732 -2760 12733 2760
rect 6811 -2761 12733 -2760
rect 6392 -2828 6488 -2812
rect 13004 -2812 13020 2812
rect 13084 -2812 13100 2812
rect 13004 -2828 13100 -2812
<< properties >>
string FIXED_BBOX 6732 -2840 12812 2840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 28.0 val 1.702k carea 2.00 cperi 0.19 nx 4 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
