magic
tech sky130A
timestamp 1730563144
<< metal1 >>
rect 100 22245 800 22275
rect 100 22105 130 22245
rect 270 22105 800 22245
rect 100 22075 800 22105
rect 700 19600 800 22075
rect 300 19400 7480 19600
rect 600 19270 7250 19300
rect 600 19130 630 19270
rect 770 19130 7250 19270
rect 600 19100 7250 19130
rect 7050 18950 7250 19100
rect 7280 18975 7480 19400
rect 8700 16270 14900 16300
rect 8700 16130 14730 16270
rect 14870 16130 14900 16270
rect 8700 16100 14900 16130
rect 7755 3810 7810 3820
rect 7755 3775 7765 3810
rect 7800 3775 7810 3810
rect 7755 3765 7810 3775
rect 7855 3810 7910 3820
rect 7855 3775 7865 3810
rect 7900 3775 7910 3810
rect 7855 3765 7910 3775
rect 7795 215 7810 3765
rect 7895 3750 7925 3765
rect 7910 285 7925 3750
rect 7910 275 11370 285
rect 7910 270 11325 275
rect 11315 240 11325 270
rect 11360 240 11370 275
rect 11315 230 11370 240
rect 7795 205 13305 215
rect 7795 200 13260 205
rect 13250 170 13260 200
rect 13295 170 13305 205
rect 13250 160 13305 170
<< via1 >>
rect 130 22105 270 22245
rect 630 19130 770 19270
rect 14730 16130 14870 16270
rect 7765 3775 7800 3810
rect 7865 3775 7900 3810
rect 11325 240 11360 275
rect 13260 170 13295 205
<< metal2 >>
rect 100 22245 300 22275
rect 100 22105 130 22245
rect 270 22105 300 22245
rect 100 22075 300 22105
rect 600 19270 800 19300
rect 600 19130 630 19270
rect 770 19130 800 19270
rect 600 19100 800 19130
rect 14700 16270 14900 16300
rect 14700 16130 14730 16270
rect 14870 16130 14900 16270
rect 14700 16100 14900 16130
rect 7755 3810 7810 3820
rect 7755 3775 7765 3810
rect 7800 3775 7810 3810
rect 7755 3765 7810 3775
rect 7855 3810 7910 3820
rect 7855 3775 7865 3810
rect 7900 3775 7910 3810
rect 7855 3765 7910 3775
rect 11315 275 11370 285
rect 11315 240 11325 275
rect 11360 240 11370 275
rect 11315 230 11370 240
rect 13250 205 13305 215
rect 13250 170 13260 205
rect 13295 170 13305 205
rect 13250 160 13305 170
<< via2 >>
rect 130 22105 270 22245
rect 630 19130 770 19270
rect 14730 16130 14870 16270
rect 7765 3775 7800 3810
rect 7865 3775 7900 3810
rect 11325 240 11360 275
rect 13260 170 13295 205
<< metal3 >>
rect 100 22245 300 22275
rect 100 22105 130 22245
rect 270 22105 300 22245
rect 100 22075 300 22105
rect 600 19270 800 19300
rect 600 19130 630 19270
rect 770 19130 800 19270
rect 600 19100 800 19130
rect 14700 16270 14900 16300
rect 14700 16130 14730 16270
rect 14870 16130 14900 16270
rect 14700 16100 14900 16130
rect 7755 3810 7810 3820
rect 7755 3775 7765 3810
rect 7800 3775 7810 3810
rect 7755 3765 7810 3775
rect 7855 3810 7910 3820
rect 7855 3775 7865 3810
rect 7900 3775 7910 3810
rect 7855 3765 7910 3775
rect 11315 275 11370 285
rect 11315 240 11325 275
rect 11360 240 11370 275
rect 11315 230 11370 240
rect 13250 205 13305 215
rect 13250 170 13260 205
rect 13295 170 13305 205
rect 13250 160 13305 170
<< via3 >>
rect 130 22105 270 22245
rect 630 19130 770 19270
rect 14730 16130 14870 16270
rect 7765 3775 7800 3810
rect 7865 3775 7900 3810
rect 11325 240 11360 275
rect 13260 170 13295 205
<< metal4 >>
rect 3067 22500 3097 22576
rect 3343 22500 3373 22576
rect 3619 22500 3649 22576
rect 3895 22500 3925 22576
rect 4171 22500 4201 22576
rect 4447 22500 4477 22576
rect 4723 22500 4753 22576
rect 4999 22500 5029 22576
rect 5275 22500 5305 22576
rect 5551 22500 5581 22576
rect 5827 22500 5857 22576
rect 6103 22500 6133 22576
rect 6379 22500 6409 22576
rect 6655 22500 6685 22576
rect 6931 22500 6961 22576
rect 7207 22500 7237 22576
rect 7483 22500 7513 22576
rect 7759 22500 7789 22576
rect 8035 22500 8065 22576
rect 8311 22500 8341 22576
rect 8587 22500 8617 22576
rect 8863 22500 8893 22576
rect 9139 22500 9169 22576
rect 9415 22500 9445 22576
rect 400 22400 9500 22500
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 100 22245 300 22275
rect 100 22105 130 22245
rect 270 22105 300 22245
rect 100 500 300 22105
rect 400 19300 600 22400
rect 400 19270 800 19300
rect 400 19130 630 19270
rect 770 19130 800 19270
rect 400 19100 800 19130
rect 400 500 600 19100
rect 14700 16270 14900 16300
rect 14700 16130 14730 16270
rect 14870 16130 14900 16270
rect 7780 3820 7810 3850
rect 7880 3820 7940 3850
rect 7755 3810 7810 3820
rect 7755 3775 7765 3810
rect 7800 3775 7810 3810
rect 7755 3765 7810 3775
rect 7855 3810 7910 3820
rect 7855 3775 7865 3810
rect 7900 3775 7910 3810
rect 7855 3765 7910 3775
rect 14700 300 14900 16130
rect 11315 275 11370 285
rect 11315 240 11325 275
rect 11360 240 11370 275
rect 11315 230 11370 240
rect 11315 100 11365 230
rect 13250 205 13305 215
rect 13250 170 13260 205
rect 13295 170 13305 205
rect 13250 100 13305 170
rect 14700 100 15300 300
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11315 90 11407 100
rect 11317 0 11407 90
rect 13249 0 13339 100
rect 15181 0 15271 100
use op_amp_3stage  op_amp_3stage_0
timestamp 1730563144
transform 1 0 22050 0 1 4195
box -20850 -3240 -7445 14825
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
rlabel metal4 400 500 600 22075 1 VGND
port 52 nsew ground bidirectional
rlabel metal4 100 500 300 22075 1 VDPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
