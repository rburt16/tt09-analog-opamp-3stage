magic
tech sky130A
magscale 1 2
timestamp 1730410385
<< pwell >>
rect -1506 -279 1506 279
<< nmos >>
rect -1310 -131 1310 69
<< ndiff >>
rect -1368 57 -1310 69
rect -1368 -119 -1356 57
rect -1322 -119 -1310 57
rect -1368 -131 -1310 -119
rect 1310 57 1368 69
rect 1310 -119 1322 57
rect 1356 -119 1368 57
rect 1310 -131 1368 -119
<< ndiffc >>
rect -1356 -119 -1322 57
rect 1322 -119 1356 57
<< psubdiff >>
rect -1470 209 1470 243
rect -1470 -209 -1436 209
rect 1436 -209 1470 209
rect -1470 -243 -1374 -209
rect 1374 -243 1470 -209
<< psubdiffcont >>
rect -1374 -243 1374 -209
<< poly >>
rect -1310 141 1310 157
rect -1310 107 -1294 141
rect 1294 107 1310 141
rect -1310 69 1310 107
rect -1310 -157 1310 -131
<< polycont >>
rect -1294 107 1294 141
<< locali >>
rect -1470 209 1470 243
rect -1470 -209 -1436 209
rect -1310 107 -1294 141
rect 1294 107 1310 141
rect -1356 57 -1322 73
rect -1356 -135 -1322 -119
rect 1322 57 1356 73
rect 1322 -135 1356 -119
rect 1436 -209 1470 209
rect -1470 -243 -1374 -209
rect 1374 -243 1470 -209
<< viali >>
rect -647 107 647 141
rect -1356 -119 -1322 57
rect 1322 -119 1356 57
rect -718 -243 718 -209
<< metal1 >>
rect -659 141 659 147
rect -659 107 -647 141
rect 647 107 659 141
rect -659 101 659 107
rect -1362 57 -1316 69
rect -1362 -119 -1356 57
rect -1322 -119 -1316 57
rect -1362 -131 -1316 -119
rect 1316 57 1362 69
rect 1316 -119 1322 57
rect 1356 -119 1362 57
rect 1316 -131 1362 -119
rect -730 -209 730 -203
rect -730 -243 -718 -209
rect 718 -243 730 -209
rect -730 -249 730 -243
<< properties >>
string FIXED_BBOX -1453 -226 1453 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 13.1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 50 viagr 0 viagl 0 viagt 0
<< end >>
