magic
tech sky130A
magscale 1 2
timestamp 1728938857
<< pwell >>
rect -4457 -510 4457 510
<< nmoslvt >>
rect -4261 -300 -3461 300
rect -3403 -300 -2603 300
rect -2545 -300 -1745 300
rect -1687 -300 -887 300
rect -829 -300 -29 300
rect 29 -300 829 300
rect 887 -300 1687 300
rect 1745 -300 2545 300
rect 2603 -300 3403 300
rect 3461 -300 4261 300
<< ndiff >>
rect -4319 288 -4261 300
rect -4319 -288 -4307 288
rect -4273 -288 -4261 288
rect -4319 -300 -4261 -288
rect -3461 288 -3403 300
rect -3461 -288 -3449 288
rect -3415 -288 -3403 288
rect -3461 -300 -3403 -288
rect -2603 288 -2545 300
rect -2603 -288 -2591 288
rect -2557 -288 -2545 288
rect -2603 -300 -2545 -288
rect -1745 288 -1687 300
rect -1745 -288 -1733 288
rect -1699 -288 -1687 288
rect -1745 -300 -1687 -288
rect -887 288 -829 300
rect -887 -288 -875 288
rect -841 -288 -829 288
rect -887 -300 -829 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 829 288 887 300
rect 829 -288 841 288
rect 875 -288 887 288
rect 829 -300 887 -288
rect 1687 288 1745 300
rect 1687 -288 1699 288
rect 1733 -288 1745 288
rect 1687 -300 1745 -288
rect 2545 288 2603 300
rect 2545 -288 2557 288
rect 2591 -288 2603 288
rect 2545 -300 2603 -288
rect 3403 288 3461 300
rect 3403 -288 3415 288
rect 3449 -288 3461 288
rect 3403 -300 3461 -288
rect 4261 288 4319 300
rect 4261 -288 4273 288
rect 4307 -288 4319 288
rect 4261 -300 4319 -288
<< ndiffc >>
rect -4307 -288 -4273 288
rect -3449 -288 -3415 288
rect -2591 -288 -2557 288
rect -1733 -288 -1699 288
rect -875 -288 -841 288
rect -17 -288 17 288
rect 841 -288 875 288
rect 1699 -288 1733 288
rect 2557 -288 2591 288
rect 3415 -288 3449 288
rect 4273 -288 4307 288
<< psubdiff >>
rect -4421 440 -4325 474
rect 4325 440 4421 474
rect -4421 378 -4387 440
rect 4387 378 4421 440
rect -4421 -440 -4387 -378
rect 4387 -440 4421 -378
rect -4421 -474 -4325 -440
rect 4325 -474 4421 -440
<< psubdiffcont >>
rect -4325 440 4325 474
rect -4421 -378 -4387 378
rect 4387 -378 4421 378
rect -4325 -474 4325 -440
<< poly >>
rect -4261 372 -3461 388
rect -4261 338 -4245 372
rect -3477 338 -3461 372
rect -4261 300 -3461 338
rect -3403 372 -2603 388
rect -3403 338 -3387 372
rect -2619 338 -2603 372
rect -3403 300 -2603 338
rect -2545 372 -1745 388
rect -2545 338 -2529 372
rect -1761 338 -1745 372
rect -2545 300 -1745 338
rect -1687 372 -887 388
rect -1687 338 -1671 372
rect -903 338 -887 372
rect -1687 300 -887 338
rect -829 372 -29 388
rect -829 338 -813 372
rect -45 338 -29 372
rect -829 300 -29 338
rect 29 372 829 388
rect 29 338 45 372
rect 813 338 829 372
rect 29 300 829 338
rect 887 372 1687 388
rect 887 338 903 372
rect 1671 338 1687 372
rect 887 300 1687 338
rect 1745 372 2545 388
rect 1745 338 1761 372
rect 2529 338 2545 372
rect 1745 300 2545 338
rect 2603 372 3403 388
rect 2603 338 2619 372
rect 3387 338 3403 372
rect 2603 300 3403 338
rect 3461 372 4261 388
rect 3461 338 3477 372
rect 4245 338 4261 372
rect 3461 300 4261 338
rect -4261 -338 -3461 -300
rect -4261 -372 -4245 -338
rect -3477 -372 -3461 -338
rect -4261 -388 -3461 -372
rect -3403 -338 -2603 -300
rect -3403 -372 -3387 -338
rect -2619 -372 -2603 -338
rect -3403 -388 -2603 -372
rect -2545 -338 -1745 -300
rect -2545 -372 -2529 -338
rect -1761 -372 -1745 -338
rect -2545 -388 -1745 -372
rect -1687 -338 -887 -300
rect -1687 -372 -1671 -338
rect -903 -372 -887 -338
rect -1687 -388 -887 -372
rect -829 -338 -29 -300
rect -829 -372 -813 -338
rect -45 -372 -29 -338
rect -829 -388 -29 -372
rect 29 -338 829 -300
rect 29 -372 45 -338
rect 813 -372 829 -338
rect 29 -388 829 -372
rect 887 -338 1687 -300
rect 887 -372 903 -338
rect 1671 -372 1687 -338
rect 887 -388 1687 -372
rect 1745 -338 2545 -300
rect 1745 -372 1761 -338
rect 2529 -372 2545 -338
rect 1745 -388 2545 -372
rect 2603 -338 3403 -300
rect 2603 -372 2619 -338
rect 3387 -372 3403 -338
rect 2603 -388 3403 -372
rect 3461 -338 4261 -300
rect 3461 -372 3477 -338
rect 4245 -372 4261 -338
rect 3461 -388 4261 -372
<< polycont >>
rect -4245 338 -3477 372
rect -3387 338 -2619 372
rect -2529 338 -1761 372
rect -1671 338 -903 372
rect -813 338 -45 372
rect 45 338 813 372
rect 903 338 1671 372
rect 1761 338 2529 372
rect 2619 338 3387 372
rect 3477 338 4245 372
rect -4245 -372 -3477 -338
rect -3387 -372 -2619 -338
rect -2529 -372 -1761 -338
rect -1671 -372 -903 -338
rect -813 -372 -45 -338
rect 45 -372 813 -338
rect 903 -372 1671 -338
rect 1761 -372 2529 -338
rect 2619 -372 3387 -338
rect 3477 -372 4245 -338
<< locali >>
rect -4421 440 -4325 474
rect 4325 440 4421 474
rect -4421 378 -4387 440
rect 4387 378 4421 440
rect -4261 338 -4245 372
rect -3477 338 -3461 372
rect -3403 338 -3387 372
rect -2619 338 -2603 372
rect -2545 338 -2529 372
rect -1761 338 -1745 372
rect -1687 338 -1671 372
rect -903 338 -887 372
rect -829 338 -813 372
rect -45 338 -29 372
rect 29 338 45 372
rect 813 338 829 372
rect 887 338 903 372
rect 1671 338 1687 372
rect 1745 338 1761 372
rect 2529 338 2545 372
rect 2603 338 2619 372
rect 3387 338 3403 372
rect 3461 338 3477 372
rect 4245 338 4261 372
rect -4307 288 -4273 304
rect -4307 -304 -4273 -288
rect -3449 288 -3415 304
rect -3449 -304 -3415 -288
rect -2591 288 -2557 304
rect -2591 -304 -2557 -288
rect -1733 288 -1699 304
rect -1733 -304 -1699 -288
rect -875 288 -841 304
rect -875 -304 -841 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 841 288 875 304
rect 841 -304 875 -288
rect 1699 288 1733 304
rect 1699 -304 1733 -288
rect 2557 288 2591 304
rect 2557 -304 2591 -288
rect 3415 288 3449 304
rect 3415 -304 3449 -288
rect 4273 288 4307 304
rect 4273 -304 4307 -288
rect -4261 -372 -4245 -338
rect -3477 -372 -3461 -338
rect -3403 -372 -3387 -338
rect -2619 -372 -2603 -338
rect -2545 -372 -2529 -338
rect -1761 -372 -1745 -338
rect -1687 -372 -1671 -338
rect -903 -372 -887 -338
rect -829 -372 -813 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 813 -372 829 -338
rect 887 -372 903 -338
rect 1671 -372 1687 -338
rect 1745 -372 1761 -338
rect 2529 -372 2545 -338
rect 2603 -372 2619 -338
rect 3387 -372 3403 -338
rect 3461 -372 3477 -338
rect 4245 -372 4261 -338
rect -4421 -440 -4387 -378
rect 4387 -440 4421 -378
rect -4421 -474 -4325 -440
rect 4325 -474 4421 -440
<< viali >>
rect -4245 338 -3477 372
rect -3387 338 -2619 372
rect -2529 338 -1761 372
rect -1671 338 -903 372
rect -813 338 -45 372
rect 45 338 813 372
rect 903 338 1671 372
rect 1761 338 2529 372
rect 2619 338 3387 372
rect 3477 338 4245 372
rect -4307 -288 -4273 288
rect -3449 -288 -3415 288
rect -2591 -288 -2557 288
rect -1733 -288 -1699 288
rect -875 -288 -841 288
rect -17 -288 17 288
rect 841 -288 875 288
rect 1699 -288 1733 288
rect 2557 -288 2591 288
rect 3415 -288 3449 288
rect 4273 -288 4307 288
rect -4245 -372 -3477 -338
rect -3387 -372 -2619 -338
rect -2529 -372 -1761 -338
rect -1671 -372 -903 -338
rect -813 -372 -45 -338
rect 45 -372 813 -338
rect 903 -372 1671 -338
rect 1761 -372 2529 -338
rect 2619 -372 3387 -338
rect 3477 -372 4245 -338
<< metal1 >>
rect -4257 372 -3465 378
rect -4257 338 -4245 372
rect -3477 338 -3465 372
rect -4257 332 -3465 338
rect -3399 372 -2607 378
rect -3399 338 -3387 372
rect -2619 338 -2607 372
rect -3399 332 -2607 338
rect -2541 372 -1749 378
rect -2541 338 -2529 372
rect -1761 338 -1749 372
rect -2541 332 -1749 338
rect -1683 372 -891 378
rect -1683 338 -1671 372
rect -903 338 -891 372
rect -1683 332 -891 338
rect -825 372 -33 378
rect -825 338 -813 372
rect -45 338 -33 372
rect -825 332 -33 338
rect 33 372 825 378
rect 33 338 45 372
rect 813 338 825 372
rect 33 332 825 338
rect 891 372 1683 378
rect 891 338 903 372
rect 1671 338 1683 372
rect 891 332 1683 338
rect 1749 372 2541 378
rect 1749 338 1761 372
rect 2529 338 2541 372
rect 1749 332 2541 338
rect 2607 372 3399 378
rect 2607 338 2619 372
rect 3387 338 3399 372
rect 2607 332 3399 338
rect 3465 372 4257 378
rect 3465 338 3477 372
rect 4245 338 4257 372
rect 3465 332 4257 338
rect -4313 288 -4267 300
rect -4313 -288 -4307 288
rect -4273 -288 -4267 288
rect -4313 -300 -4267 -288
rect -3455 288 -3409 300
rect -3455 -288 -3449 288
rect -3415 -288 -3409 288
rect -3455 -300 -3409 -288
rect -2597 288 -2551 300
rect -2597 -288 -2591 288
rect -2557 -288 -2551 288
rect -2597 -300 -2551 -288
rect -1739 288 -1693 300
rect -1739 -288 -1733 288
rect -1699 -288 -1693 288
rect -1739 -300 -1693 -288
rect -881 288 -835 300
rect -881 -288 -875 288
rect -841 -288 -835 288
rect -881 -300 -835 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 835 288 881 300
rect 835 -288 841 288
rect 875 -288 881 288
rect 835 -300 881 -288
rect 1693 288 1739 300
rect 1693 -288 1699 288
rect 1733 -288 1739 288
rect 1693 -300 1739 -288
rect 2551 288 2597 300
rect 2551 -288 2557 288
rect 2591 -288 2597 288
rect 2551 -300 2597 -288
rect 3409 288 3455 300
rect 3409 -288 3415 288
rect 3449 -288 3455 288
rect 3409 -300 3455 -288
rect 4267 288 4313 300
rect 4267 -288 4273 288
rect 4307 -288 4313 288
rect 4267 -300 4313 -288
rect -4257 -338 -3465 -332
rect -4257 -372 -4245 -338
rect -3477 -372 -3465 -338
rect -4257 -378 -3465 -372
rect -3399 -338 -2607 -332
rect -3399 -372 -3387 -338
rect -2619 -372 -2607 -338
rect -3399 -378 -2607 -372
rect -2541 -338 -1749 -332
rect -2541 -372 -2529 -338
rect -1761 -372 -1749 -338
rect -2541 -378 -1749 -372
rect -1683 -338 -891 -332
rect -1683 -372 -1671 -338
rect -903 -372 -891 -338
rect -1683 -378 -891 -372
rect -825 -338 -33 -332
rect -825 -372 -813 -338
rect -45 -372 -33 -338
rect -825 -378 -33 -372
rect 33 -338 825 -332
rect 33 -372 45 -338
rect 813 -372 825 -338
rect 33 -378 825 -372
rect 891 -338 1683 -332
rect 891 -372 903 -338
rect 1671 -372 1683 -338
rect 891 -378 1683 -372
rect 1749 -338 2541 -332
rect 1749 -372 1761 -338
rect 2529 -372 2541 -338
rect 1749 -378 2541 -372
rect 2607 -338 3399 -332
rect 2607 -372 2619 -338
rect 3387 -372 3399 -338
rect 2607 -378 3399 -372
rect 3465 -338 4257 -332
rect 3465 -372 3477 -338
rect 4245 -372 4257 -338
rect 3465 -378 4257 -372
<< properties >>
string FIXED_BBOX -4404 -457 4404 457
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3.0 l 4.0 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
