magic
tech sky130A
magscale 1 2
timestamp 1728938857
<< pwell >>
rect -596 -4191 596 4191
<< nmoslvt >>
rect -400 3381 400 3981
rect -400 2563 400 3163
rect -400 1745 400 2345
rect -400 927 400 1527
rect -400 109 400 709
rect -400 -709 400 -109
rect -400 -1527 400 -927
rect -400 -2345 400 -1745
rect -400 -3163 400 -2563
rect -400 -3981 400 -3381
<< ndiff >>
rect -458 3969 -400 3981
rect -458 3393 -446 3969
rect -412 3393 -400 3969
rect -458 3381 -400 3393
rect 400 3969 458 3981
rect 400 3393 412 3969
rect 446 3393 458 3969
rect 400 3381 458 3393
rect -458 3151 -400 3163
rect -458 2575 -446 3151
rect -412 2575 -400 3151
rect -458 2563 -400 2575
rect 400 3151 458 3163
rect 400 2575 412 3151
rect 446 2575 458 3151
rect 400 2563 458 2575
rect -458 2333 -400 2345
rect -458 1757 -446 2333
rect -412 1757 -400 2333
rect -458 1745 -400 1757
rect 400 2333 458 2345
rect 400 1757 412 2333
rect 446 1757 458 2333
rect 400 1745 458 1757
rect -458 1515 -400 1527
rect -458 939 -446 1515
rect -412 939 -400 1515
rect -458 927 -400 939
rect 400 1515 458 1527
rect 400 939 412 1515
rect 446 939 458 1515
rect 400 927 458 939
rect -458 697 -400 709
rect -458 121 -446 697
rect -412 121 -400 697
rect -458 109 -400 121
rect 400 697 458 709
rect 400 121 412 697
rect 446 121 458 697
rect 400 109 458 121
rect -458 -121 -400 -109
rect -458 -697 -446 -121
rect -412 -697 -400 -121
rect -458 -709 -400 -697
rect 400 -121 458 -109
rect 400 -697 412 -121
rect 446 -697 458 -121
rect 400 -709 458 -697
rect -458 -939 -400 -927
rect -458 -1515 -446 -939
rect -412 -1515 -400 -939
rect -458 -1527 -400 -1515
rect 400 -939 458 -927
rect 400 -1515 412 -939
rect 446 -1515 458 -939
rect 400 -1527 458 -1515
rect -458 -1757 -400 -1745
rect -458 -2333 -446 -1757
rect -412 -2333 -400 -1757
rect -458 -2345 -400 -2333
rect 400 -1757 458 -1745
rect 400 -2333 412 -1757
rect 446 -2333 458 -1757
rect 400 -2345 458 -2333
rect -458 -2575 -400 -2563
rect -458 -3151 -446 -2575
rect -412 -3151 -400 -2575
rect -458 -3163 -400 -3151
rect 400 -2575 458 -2563
rect 400 -3151 412 -2575
rect 446 -3151 458 -2575
rect 400 -3163 458 -3151
rect -458 -3393 -400 -3381
rect -458 -3969 -446 -3393
rect -412 -3969 -400 -3393
rect -458 -3981 -400 -3969
rect 400 -3393 458 -3381
rect 400 -3969 412 -3393
rect 446 -3969 458 -3393
rect 400 -3981 458 -3969
<< ndiffc >>
rect -446 3393 -412 3969
rect 412 3393 446 3969
rect -446 2575 -412 3151
rect 412 2575 446 3151
rect -446 1757 -412 2333
rect 412 1757 446 2333
rect -446 939 -412 1515
rect 412 939 446 1515
rect -446 121 -412 697
rect 412 121 446 697
rect -446 -697 -412 -121
rect 412 -697 446 -121
rect -446 -1515 -412 -939
rect 412 -1515 446 -939
rect -446 -2333 -412 -1757
rect 412 -2333 446 -1757
rect -446 -3151 -412 -2575
rect 412 -3151 446 -2575
rect -446 -3969 -412 -3393
rect 412 -3969 446 -3393
<< psubdiff >>
rect -560 4121 -464 4155
rect 464 4121 560 4155
rect -560 4059 -526 4121
rect 526 4059 560 4121
rect -560 -4121 -526 -4059
rect 526 -4121 560 -4059
rect -560 -4155 -464 -4121
rect 464 -4155 560 -4121
<< psubdiffcont >>
rect -464 4121 464 4155
rect -560 -4059 -526 4059
rect 526 -4059 560 4059
rect -464 -4155 464 -4121
<< poly >>
rect -400 4053 400 4069
rect -400 4019 -384 4053
rect 384 4019 400 4053
rect -400 3981 400 4019
rect -400 3343 400 3381
rect -400 3309 -384 3343
rect 384 3309 400 3343
rect -400 3293 400 3309
rect -400 3235 400 3251
rect -400 3201 -384 3235
rect 384 3201 400 3235
rect -400 3163 400 3201
rect -400 2525 400 2563
rect -400 2491 -384 2525
rect 384 2491 400 2525
rect -400 2475 400 2491
rect -400 2417 400 2433
rect -400 2383 -384 2417
rect 384 2383 400 2417
rect -400 2345 400 2383
rect -400 1707 400 1745
rect -400 1673 -384 1707
rect 384 1673 400 1707
rect -400 1657 400 1673
rect -400 1599 400 1615
rect -400 1565 -384 1599
rect 384 1565 400 1599
rect -400 1527 400 1565
rect -400 889 400 927
rect -400 855 -384 889
rect 384 855 400 889
rect -400 839 400 855
rect -400 781 400 797
rect -400 747 -384 781
rect 384 747 400 781
rect -400 709 400 747
rect -400 71 400 109
rect -400 37 -384 71
rect 384 37 400 71
rect -400 21 400 37
rect -400 -37 400 -21
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -400 -109 400 -71
rect -400 -747 400 -709
rect -400 -781 -384 -747
rect 384 -781 400 -747
rect -400 -797 400 -781
rect -400 -855 400 -839
rect -400 -889 -384 -855
rect 384 -889 400 -855
rect -400 -927 400 -889
rect -400 -1565 400 -1527
rect -400 -1599 -384 -1565
rect 384 -1599 400 -1565
rect -400 -1615 400 -1599
rect -400 -1673 400 -1657
rect -400 -1707 -384 -1673
rect 384 -1707 400 -1673
rect -400 -1745 400 -1707
rect -400 -2383 400 -2345
rect -400 -2417 -384 -2383
rect 384 -2417 400 -2383
rect -400 -2433 400 -2417
rect -400 -2491 400 -2475
rect -400 -2525 -384 -2491
rect 384 -2525 400 -2491
rect -400 -2563 400 -2525
rect -400 -3201 400 -3163
rect -400 -3235 -384 -3201
rect 384 -3235 400 -3201
rect -400 -3251 400 -3235
rect -400 -3309 400 -3293
rect -400 -3343 -384 -3309
rect 384 -3343 400 -3309
rect -400 -3381 400 -3343
rect -400 -4019 400 -3981
rect -400 -4053 -384 -4019
rect 384 -4053 400 -4019
rect -400 -4069 400 -4053
<< polycont >>
rect -384 4019 384 4053
rect -384 3309 384 3343
rect -384 3201 384 3235
rect -384 2491 384 2525
rect -384 2383 384 2417
rect -384 1673 384 1707
rect -384 1565 384 1599
rect -384 855 384 889
rect -384 747 384 781
rect -384 37 384 71
rect -384 -71 384 -37
rect -384 -781 384 -747
rect -384 -889 384 -855
rect -384 -1599 384 -1565
rect -384 -1707 384 -1673
rect -384 -2417 384 -2383
rect -384 -2525 384 -2491
rect -384 -3235 384 -3201
rect -384 -3343 384 -3309
rect -384 -4053 384 -4019
<< locali >>
rect -560 4121 -464 4155
rect 464 4121 560 4155
rect -560 4059 -526 4121
rect 526 4059 560 4121
rect -400 4019 -384 4053
rect 384 4019 400 4053
rect -446 3969 -412 3985
rect -446 3377 -412 3393
rect 412 3969 446 3985
rect 412 3377 446 3393
rect -400 3309 -384 3343
rect 384 3309 400 3343
rect -400 3201 -384 3235
rect 384 3201 400 3235
rect -446 3151 -412 3167
rect -446 2559 -412 2575
rect 412 3151 446 3167
rect 412 2559 446 2575
rect -400 2491 -384 2525
rect 384 2491 400 2525
rect -400 2383 -384 2417
rect 384 2383 400 2417
rect -446 2333 -412 2349
rect -446 1741 -412 1757
rect 412 2333 446 2349
rect 412 1741 446 1757
rect -400 1673 -384 1707
rect 384 1673 400 1707
rect -400 1565 -384 1599
rect 384 1565 400 1599
rect -446 1515 -412 1531
rect -446 923 -412 939
rect 412 1515 446 1531
rect 412 923 446 939
rect -400 855 -384 889
rect 384 855 400 889
rect -400 747 -384 781
rect 384 747 400 781
rect -446 697 -412 713
rect -446 105 -412 121
rect 412 697 446 713
rect 412 105 446 121
rect -400 37 -384 71
rect 384 37 400 71
rect -400 -71 -384 -37
rect 384 -71 400 -37
rect -446 -121 -412 -105
rect -446 -713 -412 -697
rect 412 -121 446 -105
rect 412 -713 446 -697
rect -400 -781 -384 -747
rect 384 -781 400 -747
rect -400 -889 -384 -855
rect 384 -889 400 -855
rect -446 -939 -412 -923
rect -446 -1531 -412 -1515
rect 412 -939 446 -923
rect 412 -1531 446 -1515
rect -400 -1599 -384 -1565
rect 384 -1599 400 -1565
rect -400 -1707 -384 -1673
rect 384 -1707 400 -1673
rect -446 -1757 -412 -1741
rect -446 -2349 -412 -2333
rect 412 -1757 446 -1741
rect 412 -2349 446 -2333
rect -400 -2417 -384 -2383
rect 384 -2417 400 -2383
rect -400 -2525 -384 -2491
rect 384 -2525 400 -2491
rect -446 -2575 -412 -2559
rect -446 -3167 -412 -3151
rect 412 -2575 446 -2559
rect 412 -3167 446 -3151
rect -400 -3235 -384 -3201
rect 384 -3235 400 -3201
rect -400 -3343 -384 -3309
rect 384 -3343 400 -3309
rect -446 -3393 -412 -3377
rect -446 -3985 -412 -3969
rect 412 -3393 446 -3377
rect 412 -3985 446 -3969
rect -400 -4053 -384 -4019
rect 384 -4053 400 -4019
rect -560 -4121 -526 -4059
rect 526 -4121 560 -4059
rect -560 -4155 -464 -4121
rect 464 -4155 560 -4121
<< viali >>
rect -384 4019 384 4053
rect -446 3393 -412 3969
rect 412 3393 446 3969
rect -384 3309 384 3343
rect -384 3201 384 3235
rect -446 2575 -412 3151
rect 412 2575 446 3151
rect -384 2491 384 2525
rect -384 2383 384 2417
rect -446 1757 -412 2333
rect 412 1757 446 2333
rect -384 1673 384 1707
rect -384 1565 384 1599
rect -446 939 -412 1515
rect 412 939 446 1515
rect -384 855 384 889
rect -384 747 384 781
rect -446 121 -412 697
rect 412 121 446 697
rect -384 37 384 71
rect -384 -71 384 -37
rect -446 -697 -412 -121
rect 412 -697 446 -121
rect -384 -781 384 -747
rect -384 -889 384 -855
rect -446 -1515 -412 -939
rect 412 -1515 446 -939
rect -384 -1599 384 -1565
rect -384 -1707 384 -1673
rect -446 -2333 -412 -1757
rect 412 -2333 446 -1757
rect -384 -2417 384 -2383
rect -384 -2525 384 -2491
rect -446 -3151 -412 -2575
rect 412 -3151 446 -2575
rect -384 -3235 384 -3201
rect -384 -3343 384 -3309
rect -446 -3969 -412 -3393
rect 412 -3969 446 -3393
rect -384 -4053 384 -4019
<< metal1 >>
rect -396 4053 396 4059
rect -396 4019 -384 4053
rect 384 4019 396 4053
rect -396 4013 396 4019
rect -452 3969 -406 3981
rect -452 3393 -446 3969
rect -412 3393 -406 3969
rect -452 3381 -406 3393
rect 406 3969 452 3981
rect 406 3393 412 3969
rect 446 3393 452 3969
rect 406 3381 452 3393
rect -396 3343 396 3349
rect -396 3309 -384 3343
rect 384 3309 396 3343
rect -396 3303 396 3309
rect -396 3235 396 3241
rect -396 3201 -384 3235
rect 384 3201 396 3235
rect -396 3195 396 3201
rect -452 3151 -406 3163
rect -452 2575 -446 3151
rect -412 2575 -406 3151
rect -452 2563 -406 2575
rect 406 3151 452 3163
rect 406 2575 412 3151
rect 446 2575 452 3151
rect 406 2563 452 2575
rect -396 2525 396 2531
rect -396 2491 -384 2525
rect 384 2491 396 2525
rect -396 2485 396 2491
rect -396 2417 396 2423
rect -396 2383 -384 2417
rect 384 2383 396 2417
rect -396 2377 396 2383
rect -452 2333 -406 2345
rect -452 1757 -446 2333
rect -412 1757 -406 2333
rect -452 1745 -406 1757
rect 406 2333 452 2345
rect 406 1757 412 2333
rect 446 1757 452 2333
rect 406 1745 452 1757
rect -396 1707 396 1713
rect -396 1673 -384 1707
rect 384 1673 396 1707
rect -396 1667 396 1673
rect -396 1599 396 1605
rect -396 1565 -384 1599
rect 384 1565 396 1599
rect -396 1559 396 1565
rect -452 1515 -406 1527
rect -452 939 -446 1515
rect -412 939 -406 1515
rect -452 927 -406 939
rect 406 1515 452 1527
rect 406 939 412 1515
rect 446 939 452 1515
rect 406 927 452 939
rect -396 889 396 895
rect -396 855 -384 889
rect 384 855 396 889
rect -396 849 396 855
rect -396 781 396 787
rect -396 747 -384 781
rect 384 747 396 781
rect -396 741 396 747
rect -452 697 -406 709
rect -452 121 -446 697
rect -412 121 -406 697
rect -452 109 -406 121
rect 406 697 452 709
rect 406 121 412 697
rect 446 121 452 697
rect 406 109 452 121
rect -396 71 396 77
rect -396 37 -384 71
rect 384 37 396 71
rect -396 31 396 37
rect -396 -37 396 -31
rect -396 -71 -384 -37
rect 384 -71 396 -37
rect -396 -77 396 -71
rect -452 -121 -406 -109
rect -452 -697 -446 -121
rect -412 -697 -406 -121
rect -452 -709 -406 -697
rect 406 -121 452 -109
rect 406 -697 412 -121
rect 446 -697 452 -121
rect 406 -709 452 -697
rect -396 -747 396 -741
rect -396 -781 -384 -747
rect 384 -781 396 -747
rect -396 -787 396 -781
rect -396 -855 396 -849
rect -396 -889 -384 -855
rect 384 -889 396 -855
rect -396 -895 396 -889
rect -452 -939 -406 -927
rect -452 -1515 -446 -939
rect -412 -1515 -406 -939
rect -452 -1527 -406 -1515
rect 406 -939 452 -927
rect 406 -1515 412 -939
rect 446 -1515 452 -939
rect 406 -1527 452 -1515
rect -396 -1565 396 -1559
rect -396 -1599 -384 -1565
rect 384 -1599 396 -1565
rect -396 -1605 396 -1599
rect -396 -1673 396 -1667
rect -396 -1707 -384 -1673
rect 384 -1707 396 -1673
rect -396 -1713 396 -1707
rect -452 -1757 -406 -1745
rect -452 -2333 -446 -1757
rect -412 -2333 -406 -1757
rect -452 -2345 -406 -2333
rect 406 -1757 452 -1745
rect 406 -2333 412 -1757
rect 446 -2333 452 -1757
rect 406 -2345 452 -2333
rect -396 -2383 396 -2377
rect -396 -2417 -384 -2383
rect 384 -2417 396 -2383
rect -396 -2423 396 -2417
rect -396 -2491 396 -2485
rect -396 -2525 -384 -2491
rect 384 -2525 396 -2491
rect -396 -2531 396 -2525
rect -452 -2575 -406 -2563
rect -452 -3151 -446 -2575
rect -412 -3151 -406 -2575
rect -452 -3163 -406 -3151
rect 406 -2575 452 -2563
rect 406 -3151 412 -2575
rect 446 -3151 452 -2575
rect 406 -3163 452 -3151
rect -396 -3201 396 -3195
rect -396 -3235 -384 -3201
rect 384 -3235 396 -3201
rect -396 -3241 396 -3235
rect -396 -3309 396 -3303
rect -396 -3343 -384 -3309
rect 384 -3343 396 -3309
rect -396 -3349 396 -3343
rect -452 -3393 -406 -3381
rect -452 -3969 -446 -3393
rect -412 -3969 -406 -3393
rect -452 -3981 -406 -3969
rect 406 -3393 452 -3381
rect 406 -3969 412 -3393
rect 446 -3969 452 -3393
rect 406 -3981 452 -3969
rect -396 -4019 396 -4013
rect -396 -4053 -384 -4019
rect 384 -4053 396 -4019
rect -396 -4059 396 -4053
<< properties >>
string FIXED_BBOX -543 -4138 543 4138
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 3.0 l 4.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
