magic
tech sky130A
magscale 1 2
timestamp 1729530615
<< error_p >>
rect -671 2199 -609 2205
rect -543 2199 -481 2205
rect -415 2199 -353 2205
rect -287 2199 -225 2205
rect -159 2199 -97 2205
rect -31 2199 31 2205
rect 97 2199 159 2205
rect 225 2199 287 2205
rect 353 2199 415 2205
rect 481 2199 543 2205
rect 609 2199 671 2205
rect -671 2165 -659 2199
rect -543 2165 -531 2199
rect -415 2165 -403 2199
rect -287 2165 -275 2199
rect -159 2165 -147 2199
rect -31 2165 -19 2199
rect 97 2165 109 2199
rect 225 2165 237 2199
rect 353 2165 365 2199
rect 481 2165 493 2199
rect 609 2165 621 2199
rect -671 2159 -609 2165
rect -543 2159 -481 2165
rect -415 2159 -353 2165
rect -287 2159 -225 2165
rect -159 2159 -97 2165
rect -31 2159 31 2165
rect 97 2159 159 2165
rect 225 2159 287 2165
rect 353 2159 415 2165
rect 481 2159 543 2165
rect 609 2159 671 2165
rect -671 71 -609 77
rect -543 71 -481 77
rect -415 71 -353 77
rect -287 71 -225 77
rect -159 71 -97 77
rect -31 71 31 77
rect 97 71 159 77
rect 225 71 287 77
rect 353 71 415 77
rect 481 71 543 77
rect 609 71 671 77
rect -671 37 -659 71
rect -543 37 -531 71
rect -415 37 -403 71
rect -287 37 -275 71
rect -159 37 -147 71
rect -31 37 -19 71
rect 97 37 109 71
rect 225 37 237 71
rect 353 37 365 71
rect 481 37 493 71
rect 609 37 621 71
rect -671 31 -609 37
rect -543 31 -481 37
rect -415 31 -353 37
rect -287 31 -225 37
rect -159 31 -97 37
rect -31 31 31 37
rect 97 31 159 37
rect 225 31 287 37
rect 353 31 415 37
rect 481 31 543 37
rect 609 31 671 37
rect -671 -37 -609 -31
rect -543 -37 -481 -31
rect -415 -37 -353 -31
rect -287 -37 -225 -31
rect -159 -37 -97 -31
rect -31 -37 31 -31
rect 97 -37 159 -31
rect 225 -37 287 -31
rect 353 -37 415 -31
rect 481 -37 543 -31
rect 609 -37 671 -31
rect -671 -71 -659 -37
rect -543 -71 -531 -37
rect -415 -71 -403 -37
rect -287 -71 -275 -37
rect -159 -71 -147 -37
rect -31 -71 -19 -37
rect 97 -71 109 -37
rect 225 -71 237 -37
rect 353 -71 365 -37
rect 481 -71 493 -37
rect 609 -71 621 -37
rect -671 -77 -609 -71
rect -543 -77 -481 -71
rect -415 -77 -353 -71
rect -287 -77 -225 -71
rect -159 -77 -97 -71
rect -31 -77 31 -71
rect 97 -77 159 -71
rect 225 -77 287 -71
rect 353 -77 415 -71
rect 481 -77 543 -71
rect 609 -77 671 -71
rect -671 -2165 -609 -2159
rect -543 -2165 -481 -2159
rect -415 -2165 -353 -2159
rect -287 -2165 -225 -2159
rect -159 -2165 -97 -2159
rect -31 -2165 31 -2159
rect 97 -2165 159 -2159
rect 225 -2165 287 -2159
rect 353 -2165 415 -2159
rect 481 -2165 543 -2159
rect 609 -2165 671 -2159
rect -671 -2199 -659 -2165
rect -543 -2199 -531 -2165
rect -415 -2199 -403 -2165
rect -287 -2199 -275 -2165
rect -159 -2199 -147 -2165
rect -31 -2199 -19 -2165
rect 97 -2199 109 -2165
rect 225 -2199 237 -2165
rect 353 -2199 365 -2165
rect 481 -2199 493 -2165
rect 609 -2199 621 -2165
rect -671 -2205 -609 -2199
rect -543 -2205 -481 -2199
rect -415 -2205 -353 -2199
rect -287 -2205 -225 -2199
rect -159 -2205 -97 -2199
rect -31 -2205 31 -2199
rect 97 -2205 159 -2199
rect 225 -2205 287 -2199
rect 353 -2205 415 -2199
rect 481 -2205 543 -2199
rect 609 -2205 671 -2199
<< nwell >>
rect -871 -2337 871 2337
<< pmoslvt >>
rect -675 118 -605 2118
rect -547 118 -477 2118
rect -419 118 -349 2118
rect -291 118 -221 2118
rect -163 118 -93 2118
rect -35 118 35 2118
rect 93 118 163 2118
rect 221 118 291 2118
rect 349 118 419 2118
rect 477 118 547 2118
rect 605 118 675 2118
rect -675 -2118 -605 -118
rect -547 -2118 -477 -118
rect -419 -2118 -349 -118
rect -291 -2118 -221 -118
rect -163 -2118 -93 -118
rect -35 -2118 35 -118
rect 93 -2118 163 -118
rect 221 -2118 291 -118
rect 349 -2118 419 -118
rect 477 -2118 547 -118
rect 605 -2118 675 -118
<< pdiff >>
rect -733 2106 -675 2118
rect -733 130 -721 2106
rect -687 130 -675 2106
rect -733 118 -675 130
rect -605 2106 -547 2118
rect -605 130 -593 2106
rect -559 130 -547 2106
rect -605 118 -547 130
rect -477 2106 -419 2118
rect -477 130 -465 2106
rect -431 130 -419 2106
rect -477 118 -419 130
rect -349 2106 -291 2118
rect -349 130 -337 2106
rect -303 130 -291 2106
rect -349 118 -291 130
rect -221 2106 -163 2118
rect -221 130 -209 2106
rect -175 130 -163 2106
rect -221 118 -163 130
rect -93 2106 -35 2118
rect -93 130 -81 2106
rect -47 130 -35 2106
rect -93 118 -35 130
rect 35 2106 93 2118
rect 35 130 47 2106
rect 81 130 93 2106
rect 35 118 93 130
rect 163 2106 221 2118
rect 163 130 175 2106
rect 209 130 221 2106
rect 163 118 221 130
rect 291 2106 349 2118
rect 291 130 303 2106
rect 337 130 349 2106
rect 291 118 349 130
rect 419 2106 477 2118
rect 419 130 431 2106
rect 465 130 477 2106
rect 419 118 477 130
rect 547 2106 605 2118
rect 547 130 559 2106
rect 593 130 605 2106
rect 547 118 605 130
rect 675 2106 733 2118
rect 675 130 687 2106
rect 721 130 733 2106
rect 675 118 733 130
rect -733 -130 -675 -118
rect -733 -2106 -721 -130
rect -687 -2106 -675 -130
rect -733 -2118 -675 -2106
rect -605 -130 -547 -118
rect -605 -2106 -593 -130
rect -559 -2106 -547 -130
rect -605 -2118 -547 -2106
rect -477 -130 -419 -118
rect -477 -2106 -465 -130
rect -431 -2106 -419 -130
rect -477 -2118 -419 -2106
rect -349 -130 -291 -118
rect -349 -2106 -337 -130
rect -303 -2106 -291 -130
rect -349 -2118 -291 -2106
rect -221 -130 -163 -118
rect -221 -2106 -209 -130
rect -175 -2106 -163 -130
rect -221 -2118 -163 -2106
rect -93 -130 -35 -118
rect -93 -2106 -81 -130
rect -47 -2106 -35 -130
rect -93 -2118 -35 -2106
rect 35 -130 93 -118
rect 35 -2106 47 -130
rect 81 -2106 93 -130
rect 35 -2118 93 -2106
rect 163 -130 221 -118
rect 163 -2106 175 -130
rect 209 -2106 221 -130
rect 163 -2118 221 -2106
rect 291 -130 349 -118
rect 291 -2106 303 -130
rect 337 -2106 349 -130
rect 291 -2118 349 -2106
rect 419 -130 477 -118
rect 419 -2106 431 -130
rect 465 -2106 477 -130
rect 419 -2118 477 -2106
rect 547 -130 605 -118
rect 547 -2106 559 -130
rect 593 -2106 605 -130
rect 547 -2118 605 -2106
rect 675 -130 733 -118
rect 675 -2106 687 -130
rect 721 -2106 733 -130
rect 675 -2118 733 -2106
<< pdiffc >>
rect -721 130 -687 2106
rect -593 130 -559 2106
rect -465 130 -431 2106
rect -337 130 -303 2106
rect -209 130 -175 2106
rect -81 130 -47 2106
rect 47 130 81 2106
rect 175 130 209 2106
rect 303 130 337 2106
rect 431 130 465 2106
rect 559 130 593 2106
rect 687 130 721 2106
rect -721 -2106 -687 -130
rect -593 -2106 -559 -130
rect -465 -2106 -431 -130
rect -337 -2106 -303 -130
rect -209 -2106 -175 -130
rect -81 -2106 -47 -130
rect 47 -2106 81 -130
rect 175 -2106 209 -130
rect 303 -2106 337 -130
rect 431 -2106 465 -130
rect 559 -2106 593 -130
rect 687 -2106 721 -130
<< nsubdiff >>
rect -835 2267 -739 2301
rect 739 2267 835 2301
rect -835 2205 -801 2267
rect 801 2205 835 2267
rect -835 -2267 -801 -2205
rect 801 -2267 835 -2205
rect -835 -2301 -739 -2267
rect 739 -2301 835 -2267
<< nsubdiffcont >>
rect -739 2267 739 2301
rect -835 -2205 -801 2205
rect 801 -2205 835 2205
rect -739 -2301 739 -2267
<< poly >>
rect -675 2199 -605 2215
rect -675 2165 -659 2199
rect -621 2165 -605 2199
rect -675 2118 -605 2165
rect -547 2199 -477 2215
rect -547 2165 -531 2199
rect -493 2165 -477 2199
rect -547 2118 -477 2165
rect -419 2199 -349 2215
rect -419 2165 -403 2199
rect -365 2165 -349 2199
rect -419 2118 -349 2165
rect -291 2199 -221 2215
rect -291 2165 -275 2199
rect -237 2165 -221 2199
rect -291 2118 -221 2165
rect -163 2199 -93 2215
rect -163 2165 -147 2199
rect -109 2165 -93 2199
rect -163 2118 -93 2165
rect -35 2199 35 2215
rect -35 2165 -19 2199
rect 19 2165 35 2199
rect -35 2118 35 2165
rect 93 2199 163 2215
rect 93 2165 109 2199
rect 147 2165 163 2199
rect 93 2118 163 2165
rect 221 2199 291 2215
rect 221 2165 237 2199
rect 275 2165 291 2199
rect 221 2118 291 2165
rect 349 2199 419 2215
rect 349 2165 365 2199
rect 403 2165 419 2199
rect 349 2118 419 2165
rect 477 2199 547 2215
rect 477 2165 493 2199
rect 531 2165 547 2199
rect 477 2118 547 2165
rect 605 2199 675 2215
rect 605 2165 621 2199
rect 659 2165 675 2199
rect 605 2118 675 2165
rect -675 71 -605 118
rect -675 37 -659 71
rect -621 37 -605 71
rect -675 21 -605 37
rect -547 71 -477 118
rect -547 37 -531 71
rect -493 37 -477 71
rect -547 21 -477 37
rect -419 71 -349 118
rect -419 37 -403 71
rect -365 37 -349 71
rect -419 21 -349 37
rect -291 71 -221 118
rect -291 37 -275 71
rect -237 37 -221 71
rect -291 21 -221 37
rect -163 71 -93 118
rect -163 37 -147 71
rect -109 37 -93 71
rect -163 21 -93 37
rect -35 71 35 118
rect -35 37 -19 71
rect 19 37 35 71
rect -35 21 35 37
rect 93 71 163 118
rect 93 37 109 71
rect 147 37 163 71
rect 93 21 163 37
rect 221 71 291 118
rect 221 37 237 71
rect 275 37 291 71
rect 221 21 291 37
rect 349 71 419 118
rect 349 37 365 71
rect 403 37 419 71
rect 349 21 419 37
rect 477 71 547 118
rect 477 37 493 71
rect 531 37 547 71
rect 477 21 547 37
rect 605 71 675 118
rect 605 37 621 71
rect 659 37 675 71
rect 605 21 675 37
rect -675 -37 -605 -21
rect -675 -71 -659 -37
rect -621 -71 -605 -37
rect -675 -118 -605 -71
rect -547 -37 -477 -21
rect -547 -71 -531 -37
rect -493 -71 -477 -37
rect -547 -118 -477 -71
rect -419 -37 -349 -21
rect -419 -71 -403 -37
rect -365 -71 -349 -37
rect -419 -118 -349 -71
rect -291 -37 -221 -21
rect -291 -71 -275 -37
rect -237 -71 -221 -37
rect -291 -118 -221 -71
rect -163 -37 -93 -21
rect -163 -71 -147 -37
rect -109 -71 -93 -37
rect -163 -118 -93 -71
rect -35 -37 35 -21
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -35 -118 35 -71
rect 93 -37 163 -21
rect 93 -71 109 -37
rect 147 -71 163 -37
rect 93 -118 163 -71
rect 221 -37 291 -21
rect 221 -71 237 -37
rect 275 -71 291 -37
rect 221 -118 291 -71
rect 349 -37 419 -21
rect 349 -71 365 -37
rect 403 -71 419 -37
rect 349 -118 419 -71
rect 477 -37 547 -21
rect 477 -71 493 -37
rect 531 -71 547 -37
rect 477 -118 547 -71
rect 605 -37 675 -21
rect 605 -71 621 -37
rect 659 -71 675 -37
rect 605 -118 675 -71
rect -675 -2165 -605 -2118
rect -675 -2199 -659 -2165
rect -621 -2199 -605 -2165
rect -675 -2215 -605 -2199
rect -547 -2165 -477 -2118
rect -547 -2199 -531 -2165
rect -493 -2199 -477 -2165
rect -547 -2215 -477 -2199
rect -419 -2165 -349 -2118
rect -419 -2199 -403 -2165
rect -365 -2199 -349 -2165
rect -419 -2215 -349 -2199
rect -291 -2165 -221 -2118
rect -291 -2199 -275 -2165
rect -237 -2199 -221 -2165
rect -291 -2215 -221 -2199
rect -163 -2165 -93 -2118
rect -163 -2199 -147 -2165
rect -109 -2199 -93 -2165
rect -163 -2215 -93 -2199
rect -35 -2165 35 -2118
rect -35 -2199 -19 -2165
rect 19 -2199 35 -2165
rect -35 -2215 35 -2199
rect 93 -2165 163 -2118
rect 93 -2199 109 -2165
rect 147 -2199 163 -2165
rect 93 -2215 163 -2199
rect 221 -2165 291 -2118
rect 221 -2199 237 -2165
rect 275 -2199 291 -2165
rect 221 -2215 291 -2199
rect 349 -2165 419 -2118
rect 349 -2199 365 -2165
rect 403 -2199 419 -2165
rect 349 -2215 419 -2199
rect 477 -2165 547 -2118
rect 477 -2199 493 -2165
rect 531 -2199 547 -2165
rect 477 -2215 547 -2199
rect 605 -2165 675 -2118
rect 605 -2199 621 -2165
rect 659 -2199 675 -2165
rect 605 -2215 675 -2199
<< polycont >>
rect -659 2165 -621 2199
rect -531 2165 -493 2199
rect -403 2165 -365 2199
rect -275 2165 -237 2199
rect -147 2165 -109 2199
rect -19 2165 19 2199
rect 109 2165 147 2199
rect 237 2165 275 2199
rect 365 2165 403 2199
rect 493 2165 531 2199
rect 621 2165 659 2199
rect -659 37 -621 71
rect -531 37 -493 71
rect -403 37 -365 71
rect -275 37 -237 71
rect -147 37 -109 71
rect -19 37 19 71
rect 109 37 147 71
rect 237 37 275 71
rect 365 37 403 71
rect 493 37 531 71
rect 621 37 659 71
rect -659 -71 -621 -37
rect -531 -71 -493 -37
rect -403 -71 -365 -37
rect -275 -71 -237 -37
rect -147 -71 -109 -37
rect -19 -71 19 -37
rect 109 -71 147 -37
rect 237 -71 275 -37
rect 365 -71 403 -37
rect 493 -71 531 -37
rect 621 -71 659 -37
rect -659 -2199 -621 -2165
rect -531 -2199 -493 -2165
rect -403 -2199 -365 -2165
rect -275 -2199 -237 -2165
rect -147 -2199 -109 -2165
rect -19 -2199 19 -2165
rect 109 -2199 147 -2165
rect 237 -2199 275 -2165
rect 365 -2199 403 -2165
rect 493 -2199 531 -2165
rect 621 -2199 659 -2165
<< locali >>
rect -835 2267 -739 2301
rect 739 2267 835 2301
rect -835 2205 -801 2267
rect 801 2205 835 2267
rect -675 2165 -659 2199
rect -621 2165 -605 2199
rect -547 2165 -531 2199
rect -493 2165 -477 2199
rect -419 2165 -403 2199
rect -365 2165 -349 2199
rect -291 2165 -275 2199
rect -237 2165 -221 2199
rect -163 2165 -147 2199
rect -109 2165 -93 2199
rect -35 2165 -19 2199
rect 19 2165 35 2199
rect 93 2165 109 2199
rect 147 2165 163 2199
rect 221 2165 237 2199
rect 275 2165 291 2199
rect 349 2165 365 2199
rect 403 2165 419 2199
rect 477 2165 493 2199
rect 531 2165 547 2199
rect 605 2165 621 2199
rect 659 2165 675 2199
rect -721 2106 -687 2122
rect -721 114 -687 130
rect -593 2106 -559 2122
rect -593 114 -559 130
rect -465 2106 -431 2122
rect -465 114 -431 130
rect -337 2106 -303 2122
rect -337 114 -303 130
rect -209 2106 -175 2122
rect -209 114 -175 130
rect -81 2106 -47 2122
rect -81 114 -47 130
rect 47 2106 81 2122
rect 47 114 81 130
rect 175 2106 209 2122
rect 175 114 209 130
rect 303 2106 337 2122
rect 303 114 337 130
rect 431 2106 465 2122
rect 431 114 465 130
rect 559 2106 593 2122
rect 559 114 593 130
rect 687 2106 721 2122
rect 687 114 721 130
rect -675 37 -659 71
rect -621 37 -605 71
rect -547 37 -531 71
rect -493 37 -477 71
rect -419 37 -403 71
rect -365 37 -349 71
rect -291 37 -275 71
rect -237 37 -221 71
rect -163 37 -147 71
rect -109 37 -93 71
rect -35 37 -19 71
rect 19 37 35 71
rect 93 37 109 71
rect 147 37 163 71
rect 221 37 237 71
rect 275 37 291 71
rect 349 37 365 71
rect 403 37 419 71
rect 477 37 493 71
rect 531 37 547 71
rect 605 37 621 71
rect 659 37 675 71
rect -675 -71 -659 -37
rect -621 -71 -605 -37
rect -547 -71 -531 -37
rect -493 -71 -477 -37
rect -419 -71 -403 -37
rect -365 -71 -349 -37
rect -291 -71 -275 -37
rect -237 -71 -221 -37
rect -163 -71 -147 -37
rect -109 -71 -93 -37
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect 93 -71 109 -37
rect 147 -71 163 -37
rect 221 -71 237 -37
rect 275 -71 291 -37
rect 349 -71 365 -37
rect 403 -71 419 -37
rect 477 -71 493 -37
rect 531 -71 547 -37
rect 605 -71 621 -37
rect 659 -71 675 -37
rect -721 -130 -687 -114
rect -721 -2122 -687 -2106
rect -593 -130 -559 -114
rect -593 -2122 -559 -2106
rect -465 -130 -431 -114
rect -465 -2122 -431 -2106
rect -337 -130 -303 -114
rect -337 -2122 -303 -2106
rect -209 -130 -175 -114
rect -209 -2122 -175 -2106
rect -81 -130 -47 -114
rect -81 -2122 -47 -2106
rect 47 -130 81 -114
rect 47 -2122 81 -2106
rect 175 -130 209 -114
rect 175 -2122 209 -2106
rect 303 -130 337 -114
rect 303 -2122 337 -2106
rect 431 -130 465 -114
rect 431 -2122 465 -2106
rect 559 -130 593 -114
rect 559 -2122 593 -2106
rect 687 -130 721 -114
rect 687 -2122 721 -2106
rect -675 -2199 -659 -2165
rect -621 -2199 -605 -2165
rect -547 -2199 -531 -2165
rect -493 -2199 -477 -2165
rect -419 -2199 -403 -2165
rect -365 -2199 -349 -2165
rect -291 -2199 -275 -2165
rect -237 -2199 -221 -2165
rect -163 -2199 -147 -2165
rect -109 -2199 -93 -2165
rect -35 -2199 -19 -2165
rect 19 -2199 35 -2165
rect 93 -2199 109 -2165
rect 147 -2199 163 -2165
rect 221 -2199 237 -2165
rect 275 -2199 291 -2165
rect 349 -2199 365 -2165
rect 403 -2199 419 -2165
rect 477 -2199 493 -2165
rect 531 -2199 547 -2165
rect 605 -2199 621 -2165
rect 659 -2199 675 -2165
rect -835 -2267 -801 -2205
rect 801 -2267 835 -2205
rect -835 -2301 -739 -2267
rect 739 -2301 835 -2267
<< viali >>
rect -659 2165 -621 2199
rect -531 2165 -493 2199
rect -403 2165 -365 2199
rect -275 2165 -237 2199
rect -147 2165 -109 2199
rect -19 2165 19 2199
rect 109 2165 147 2199
rect 237 2165 275 2199
rect 365 2165 403 2199
rect 493 2165 531 2199
rect 621 2165 659 2199
rect -721 130 -687 2106
rect -593 130 -559 2106
rect -465 130 -431 2106
rect -337 130 -303 2106
rect -209 130 -175 2106
rect -81 130 -47 2106
rect 47 130 81 2106
rect 175 130 209 2106
rect 303 130 337 2106
rect 431 130 465 2106
rect 559 130 593 2106
rect 687 130 721 2106
rect -659 37 -621 71
rect -531 37 -493 71
rect -403 37 -365 71
rect -275 37 -237 71
rect -147 37 -109 71
rect -19 37 19 71
rect 109 37 147 71
rect 237 37 275 71
rect 365 37 403 71
rect 493 37 531 71
rect 621 37 659 71
rect -659 -71 -621 -37
rect -531 -71 -493 -37
rect -403 -71 -365 -37
rect -275 -71 -237 -37
rect -147 -71 -109 -37
rect -19 -71 19 -37
rect 109 -71 147 -37
rect 237 -71 275 -37
rect 365 -71 403 -37
rect 493 -71 531 -37
rect 621 -71 659 -37
rect -721 -2106 -687 -130
rect -593 -2106 -559 -130
rect -465 -2106 -431 -130
rect -337 -2106 -303 -130
rect -209 -2106 -175 -130
rect -81 -2106 -47 -130
rect 47 -2106 81 -130
rect 175 -2106 209 -130
rect 303 -2106 337 -130
rect 431 -2106 465 -130
rect 559 -2106 593 -130
rect 687 -2106 721 -130
rect -659 -2199 -621 -2165
rect -531 -2199 -493 -2165
rect -403 -2199 -365 -2165
rect -275 -2199 -237 -2165
rect -147 -2199 -109 -2165
rect -19 -2199 19 -2165
rect 109 -2199 147 -2165
rect 237 -2199 275 -2165
rect 365 -2199 403 -2165
rect 493 -2199 531 -2165
rect 621 -2199 659 -2165
<< metal1 >>
rect -671 2199 -609 2205
rect -671 2165 -659 2199
rect -621 2165 -609 2199
rect -671 2159 -609 2165
rect -543 2199 -481 2205
rect -543 2165 -531 2199
rect -493 2165 -481 2199
rect -543 2159 -481 2165
rect -415 2199 -353 2205
rect -415 2165 -403 2199
rect -365 2165 -353 2199
rect -415 2159 -353 2165
rect -287 2199 -225 2205
rect -287 2165 -275 2199
rect -237 2165 -225 2199
rect -287 2159 -225 2165
rect -159 2199 -97 2205
rect -159 2165 -147 2199
rect -109 2165 -97 2199
rect -159 2159 -97 2165
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect 19 2165 31 2199
rect -31 2159 31 2165
rect 97 2199 159 2205
rect 97 2165 109 2199
rect 147 2165 159 2199
rect 97 2159 159 2165
rect 225 2199 287 2205
rect 225 2165 237 2199
rect 275 2165 287 2199
rect 225 2159 287 2165
rect 353 2199 415 2205
rect 353 2165 365 2199
rect 403 2165 415 2199
rect 353 2159 415 2165
rect 481 2199 543 2205
rect 481 2165 493 2199
rect 531 2165 543 2199
rect 481 2159 543 2165
rect 609 2199 671 2205
rect 609 2165 621 2199
rect 659 2165 671 2199
rect 609 2159 671 2165
rect -727 2106 -681 2118
rect -727 130 -721 2106
rect -687 130 -681 2106
rect -727 118 -681 130
rect -599 2106 -553 2118
rect -599 130 -593 2106
rect -559 130 -553 2106
rect -599 118 -553 130
rect -471 2106 -425 2118
rect -471 130 -465 2106
rect -431 130 -425 2106
rect -471 118 -425 130
rect -343 2106 -297 2118
rect -343 130 -337 2106
rect -303 130 -297 2106
rect -343 118 -297 130
rect -215 2106 -169 2118
rect -215 130 -209 2106
rect -175 130 -169 2106
rect -215 118 -169 130
rect -87 2106 -41 2118
rect -87 130 -81 2106
rect -47 130 -41 2106
rect -87 118 -41 130
rect 41 2106 87 2118
rect 41 130 47 2106
rect 81 130 87 2106
rect 41 118 87 130
rect 169 2106 215 2118
rect 169 130 175 2106
rect 209 130 215 2106
rect 169 118 215 130
rect 297 2106 343 2118
rect 297 130 303 2106
rect 337 130 343 2106
rect 297 118 343 130
rect 425 2106 471 2118
rect 425 130 431 2106
rect 465 130 471 2106
rect 425 118 471 130
rect 553 2106 599 2118
rect 553 130 559 2106
rect 593 130 599 2106
rect 553 118 599 130
rect 681 2106 727 2118
rect 681 130 687 2106
rect 721 130 727 2106
rect 681 118 727 130
rect -671 71 -609 77
rect -671 37 -659 71
rect -621 37 -609 71
rect -671 31 -609 37
rect -543 71 -481 77
rect -543 37 -531 71
rect -493 37 -481 71
rect -543 31 -481 37
rect -415 71 -353 77
rect -415 37 -403 71
rect -365 37 -353 71
rect -415 31 -353 37
rect -287 71 -225 77
rect -287 37 -275 71
rect -237 37 -225 71
rect -287 31 -225 37
rect -159 71 -97 77
rect -159 37 -147 71
rect -109 37 -97 71
rect -159 31 -97 37
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect 97 71 159 77
rect 97 37 109 71
rect 147 37 159 71
rect 97 31 159 37
rect 225 71 287 77
rect 225 37 237 71
rect 275 37 287 71
rect 225 31 287 37
rect 353 71 415 77
rect 353 37 365 71
rect 403 37 415 71
rect 353 31 415 37
rect 481 71 543 77
rect 481 37 493 71
rect 531 37 543 71
rect 481 31 543 37
rect 609 71 671 77
rect 609 37 621 71
rect 659 37 671 71
rect 609 31 671 37
rect -671 -37 -609 -31
rect -671 -71 -659 -37
rect -621 -71 -609 -37
rect -671 -77 -609 -71
rect -543 -37 -481 -31
rect -543 -71 -531 -37
rect -493 -71 -481 -37
rect -543 -77 -481 -71
rect -415 -37 -353 -31
rect -415 -71 -403 -37
rect -365 -71 -353 -37
rect -415 -77 -353 -71
rect -287 -37 -225 -31
rect -287 -71 -275 -37
rect -237 -71 -225 -37
rect -287 -77 -225 -71
rect -159 -37 -97 -31
rect -159 -71 -147 -37
rect -109 -71 -97 -37
rect -159 -77 -97 -71
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect 97 -37 159 -31
rect 97 -71 109 -37
rect 147 -71 159 -37
rect 97 -77 159 -71
rect 225 -37 287 -31
rect 225 -71 237 -37
rect 275 -71 287 -37
rect 225 -77 287 -71
rect 353 -37 415 -31
rect 353 -71 365 -37
rect 403 -71 415 -37
rect 353 -77 415 -71
rect 481 -37 543 -31
rect 481 -71 493 -37
rect 531 -71 543 -37
rect 481 -77 543 -71
rect 609 -37 671 -31
rect 609 -71 621 -37
rect 659 -71 671 -37
rect 609 -77 671 -71
rect -727 -130 -681 -118
rect -727 -2106 -721 -130
rect -687 -2106 -681 -130
rect -727 -2118 -681 -2106
rect -599 -130 -553 -118
rect -599 -2106 -593 -130
rect -559 -2106 -553 -130
rect -599 -2118 -553 -2106
rect -471 -130 -425 -118
rect -471 -2106 -465 -130
rect -431 -2106 -425 -130
rect -471 -2118 -425 -2106
rect -343 -130 -297 -118
rect -343 -2106 -337 -130
rect -303 -2106 -297 -130
rect -343 -2118 -297 -2106
rect -215 -130 -169 -118
rect -215 -2106 -209 -130
rect -175 -2106 -169 -130
rect -215 -2118 -169 -2106
rect -87 -130 -41 -118
rect -87 -2106 -81 -130
rect -47 -2106 -41 -130
rect -87 -2118 -41 -2106
rect 41 -130 87 -118
rect 41 -2106 47 -130
rect 81 -2106 87 -130
rect 41 -2118 87 -2106
rect 169 -130 215 -118
rect 169 -2106 175 -130
rect 209 -2106 215 -130
rect 169 -2118 215 -2106
rect 297 -130 343 -118
rect 297 -2106 303 -130
rect 337 -2106 343 -130
rect 297 -2118 343 -2106
rect 425 -130 471 -118
rect 425 -2106 431 -130
rect 465 -2106 471 -130
rect 425 -2118 471 -2106
rect 553 -130 599 -118
rect 553 -2106 559 -130
rect 593 -2106 599 -130
rect 553 -2118 599 -2106
rect 681 -130 727 -118
rect 681 -2106 687 -130
rect 721 -2106 727 -130
rect 681 -2118 727 -2106
rect -671 -2165 -609 -2159
rect -671 -2199 -659 -2165
rect -621 -2199 -609 -2165
rect -671 -2205 -609 -2199
rect -543 -2165 -481 -2159
rect -543 -2199 -531 -2165
rect -493 -2199 -481 -2165
rect -543 -2205 -481 -2199
rect -415 -2165 -353 -2159
rect -415 -2199 -403 -2165
rect -365 -2199 -353 -2165
rect -415 -2205 -353 -2199
rect -287 -2165 -225 -2159
rect -287 -2199 -275 -2165
rect -237 -2199 -225 -2165
rect -287 -2205 -225 -2199
rect -159 -2165 -97 -2159
rect -159 -2199 -147 -2165
rect -109 -2199 -97 -2165
rect -159 -2205 -97 -2199
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect 19 -2199 31 -2165
rect -31 -2205 31 -2199
rect 97 -2165 159 -2159
rect 97 -2199 109 -2165
rect 147 -2199 159 -2165
rect 97 -2205 159 -2199
rect 225 -2165 287 -2159
rect 225 -2199 237 -2165
rect 275 -2199 287 -2165
rect 225 -2205 287 -2199
rect 353 -2165 415 -2159
rect 353 -2199 365 -2165
rect 403 -2199 415 -2165
rect 353 -2205 415 -2199
rect 481 -2165 543 -2159
rect 481 -2199 493 -2165
rect 531 -2199 543 -2165
rect 481 -2205 543 -2199
rect 609 -2165 671 -2159
rect 609 -2199 621 -2165
rect 659 -2199 671 -2165
rect 609 -2205 671 -2199
<< properties >>
string FIXED_BBOX -818 -2284 818 2284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 2 nf 11 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
