magic
tech sky130A
magscale 1 2
timestamp 1730569394
<< nwell >>
rect -3335 -2219 3335 2219
<< pmoslvt >>
rect -3139 -2000 -2999 2000
rect -2941 -2000 -2801 2000
rect -2743 -2000 -2603 2000
rect -2545 -2000 -2405 2000
rect -2347 -2000 -2207 2000
rect -2149 -2000 -2009 2000
rect -1951 -2000 -1811 2000
rect -1753 -2000 -1613 2000
rect -1555 -2000 -1415 2000
rect -1357 -2000 -1217 2000
rect -1159 -2000 -1019 2000
rect -961 -2000 -821 2000
rect -763 -2000 -623 2000
rect -565 -2000 -425 2000
rect -367 -2000 -227 2000
rect -169 -2000 -29 2000
rect 29 -2000 169 2000
rect 227 -2000 367 2000
rect 425 -2000 565 2000
rect 623 -2000 763 2000
rect 821 -2000 961 2000
rect 1019 -2000 1159 2000
rect 1217 -2000 1357 2000
rect 1415 -2000 1555 2000
rect 1613 -2000 1753 2000
rect 1811 -2000 1951 2000
rect 2009 -2000 2149 2000
rect 2207 -2000 2347 2000
rect 2405 -2000 2545 2000
rect 2603 -2000 2743 2000
rect 2801 -2000 2941 2000
rect 2999 -2000 3139 2000
<< pdiff >>
rect -3197 1392 -3139 2000
rect -3197 -1392 -3185 1392
rect -3151 -1392 -3139 1392
rect -3197 -2000 -3139 -1392
rect -2999 1392 -2941 2000
rect -2999 -1392 -2987 1392
rect -2953 -1392 -2941 1392
rect -2999 -2000 -2941 -1392
rect -2801 1392 -2743 2000
rect -2801 -1392 -2789 1392
rect -2755 -1392 -2743 1392
rect -2801 -2000 -2743 -1392
rect -2603 1392 -2545 2000
rect -2603 -1392 -2591 1392
rect -2557 -1392 -2545 1392
rect -2603 -2000 -2545 -1392
rect -2405 1392 -2347 2000
rect -2405 -1392 -2393 1392
rect -2359 -1392 -2347 1392
rect -2405 -2000 -2347 -1392
rect -2207 1392 -2149 2000
rect -2207 -1392 -2195 1392
rect -2161 -1392 -2149 1392
rect -2207 -2000 -2149 -1392
rect -2009 1392 -1951 2000
rect -2009 -1392 -1997 1392
rect -1963 -1392 -1951 1392
rect -2009 -2000 -1951 -1392
rect -1811 1392 -1753 2000
rect -1811 -1392 -1799 1392
rect -1765 -1392 -1753 1392
rect -1811 -2000 -1753 -1392
rect -1613 1392 -1555 2000
rect -1613 -1392 -1601 1392
rect -1567 -1392 -1555 1392
rect -1613 -2000 -1555 -1392
rect -1415 1392 -1357 2000
rect -1415 -1392 -1403 1392
rect -1369 -1392 -1357 1392
rect -1415 -2000 -1357 -1392
rect -1217 1392 -1159 2000
rect -1217 -1392 -1205 1392
rect -1171 -1392 -1159 1392
rect -1217 -2000 -1159 -1392
rect -1019 1392 -961 2000
rect -1019 -1392 -1007 1392
rect -973 -1392 -961 1392
rect -1019 -2000 -961 -1392
rect -821 1392 -763 2000
rect -821 -1392 -809 1392
rect -775 -1392 -763 1392
rect -821 -2000 -763 -1392
rect -623 1392 -565 2000
rect -623 -1392 -611 1392
rect -577 -1392 -565 1392
rect -623 -2000 -565 -1392
rect -425 1392 -367 2000
rect -425 -1392 -413 1392
rect -379 -1392 -367 1392
rect -425 -2000 -367 -1392
rect -227 1392 -169 2000
rect -227 -1392 -215 1392
rect -181 -1392 -169 1392
rect -227 -2000 -169 -1392
rect -29 1392 29 2000
rect -29 -1392 -17 1392
rect 17 -1392 29 1392
rect -29 -2000 29 -1392
rect 169 1392 227 2000
rect 169 -1392 181 1392
rect 215 -1392 227 1392
rect 169 -2000 227 -1392
rect 367 1392 425 2000
rect 367 -1392 379 1392
rect 413 -1392 425 1392
rect 367 -2000 425 -1392
rect 565 1392 623 2000
rect 565 -1392 577 1392
rect 611 -1392 623 1392
rect 565 -2000 623 -1392
rect 763 1392 821 2000
rect 763 -1392 775 1392
rect 809 -1392 821 1392
rect 763 -2000 821 -1392
rect 961 1392 1019 2000
rect 961 -1392 973 1392
rect 1007 -1392 1019 1392
rect 961 -2000 1019 -1392
rect 1159 1392 1217 2000
rect 1159 -1392 1171 1392
rect 1205 -1392 1217 1392
rect 1159 -2000 1217 -1392
rect 1357 1392 1415 2000
rect 1357 -1392 1369 1392
rect 1403 -1392 1415 1392
rect 1357 -2000 1415 -1392
rect 1555 1392 1613 2000
rect 1555 -1392 1567 1392
rect 1601 -1392 1613 1392
rect 1555 -2000 1613 -1392
rect 1753 1392 1811 2000
rect 1753 -1392 1765 1392
rect 1799 -1392 1811 1392
rect 1753 -2000 1811 -1392
rect 1951 1392 2009 2000
rect 1951 -1392 1963 1392
rect 1997 -1392 2009 1392
rect 1951 -2000 2009 -1392
rect 2149 1392 2207 2000
rect 2149 -1392 2161 1392
rect 2195 -1392 2207 1392
rect 2149 -2000 2207 -1392
rect 2347 1392 2405 2000
rect 2347 -1392 2359 1392
rect 2393 -1392 2405 1392
rect 2347 -2000 2405 -1392
rect 2545 1392 2603 2000
rect 2545 -1392 2557 1392
rect 2591 -1392 2603 1392
rect 2545 -2000 2603 -1392
rect 2743 1392 2801 2000
rect 2743 -1392 2755 1392
rect 2789 -1392 2801 1392
rect 2743 -2000 2801 -1392
rect 2941 1392 2999 2000
rect 2941 -1392 2953 1392
rect 2987 -1392 2999 1392
rect 2941 -2000 2999 -1392
rect 3139 1392 3197 2000
rect 3139 -1392 3151 1392
rect 3185 -1392 3197 1392
rect 3139 -2000 3197 -1392
<< pdiffc >>
rect -3185 -1392 -3151 1392
rect -2987 -1392 -2953 1392
rect -2789 -1392 -2755 1392
rect -2591 -1392 -2557 1392
rect -2393 -1392 -2359 1392
rect -2195 -1392 -2161 1392
rect -1997 -1392 -1963 1392
rect -1799 -1392 -1765 1392
rect -1601 -1392 -1567 1392
rect -1403 -1392 -1369 1392
rect -1205 -1392 -1171 1392
rect -1007 -1392 -973 1392
rect -809 -1392 -775 1392
rect -611 -1392 -577 1392
rect -413 -1392 -379 1392
rect -215 -1392 -181 1392
rect -17 -1392 17 1392
rect 181 -1392 215 1392
rect 379 -1392 413 1392
rect 577 -1392 611 1392
rect 775 -1392 809 1392
rect 973 -1392 1007 1392
rect 1171 -1392 1205 1392
rect 1369 -1392 1403 1392
rect 1567 -1392 1601 1392
rect 1765 -1392 1799 1392
rect 1963 -1392 1997 1392
rect 2161 -1392 2195 1392
rect 2359 -1392 2393 1392
rect 2557 -1392 2591 1392
rect 2755 -1392 2789 1392
rect 2953 -1392 2987 1392
rect 3151 -1392 3185 1392
<< nsubdiff >>
rect -3299 2149 -2242 2183
rect 2242 2149 3299 2183
rect -3299 1461 -3265 2149
rect -3299 -2149 -3265 -1461
rect 3265 1461 3299 2149
rect 3265 -2149 3299 -1461
rect -3299 -2183 -2242 -2149
rect 2242 -2183 3299 -2149
<< nsubdiffcont >>
rect -2242 2149 2242 2183
rect -3299 -1461 -3265 1461
rect 3265 -1461 3299 1461
rect -2242 -2183 2242 -2149
<< poly >>
rect -3123 2081 -3015 2097
rect -3123 2064 -3107 2081
rect -3139 2047 -3107 2064
rect -3031 2064 -3015 2081
rect -2925 2081 -2817 2097
rect -2925 2064 -2909 2081
rect -3031 2047 -2999 2064
rect -3139 2000 -2999 2047
rect -2941 2047 -2909 2064
rect -2833 2064 -2817 2081
rect -2727 2081 -2619 2097
rect -2727 2064 -2711 2081
rect -2833 2047 -2801 2064
rect -2941 2000 -2801 2047
rect -2743 2047 -2711 2064
rect -2635 2064 -2619 2081
rect -2529 2081 -2421 2097
rect -2529 2064 -2513 2081
rect -2635 2047 -2603 2064
rect -2743 2000 -2603 2047
rect -2545 2047 -2513 2064
rect -2437 2064 -2421 2081
rect -2331 2081 -2223 2097
rect -2331 2064 -2315 2081
rect -2437 2047 -2405 2064
rect -2545 2000 -2405 2047
rect -2347 2047 -2315 2064
rect -2239 2064 -2223 2081
rect -2133 2081 -2025 2097
rect -2133 2064 -2117 2081
rect -2239 2047 -2207 2064
rect -2347 2000 -2207 2047
rect -2149 2047 -2117 2064
rect -2041 2064 -2025 2081
rect -1935 2081 -1827 2097
rect -1935 2064 -1919 2081
rect -2041 2047 -2009 2064
rect -2149 2000 -2009 2047
rect -1951 2047 -1919 2064
rect -1843 2064 -1827 2081
rect -1737 2081 -1629 2097
rect -1737 2064 -1721 2081
rect -1843 2047 -1811 2064
rect -1951 2000 -1811 2047
rect -1753 2047 -1721 2064
rect -1645 2064 -1629 2081
rect -1539 2081 -1431 2097
rect -1539 2064 -1523 2081
rect -1645 2047 -1613 2064
rect -1753 2000 -1613 2047
rect -1555 2047 -1523 2064
rect -1447 2064 -1431 2081
rect -1341 2081 -1233 2097
rect -1341 2064 -1325 2081
rect -1447 2047 -1415 2064
rect -1555 2000 -1415 2047
rect -1357 2047 -1325 2064
rect -1249 2064 -1233 2081
rect -1143 2081 -1035 2097
rect -1143 2064 -1127 2081
rect -1249 2047 -1217 2064
rect -1357 2000 -1217 2047
rect -1159 2047 -1127 2064
rect -1051 2064 -1035 2081
rect -945 2081 -837 2097
rect -945 2064 -929 2081
rect -1051 2047 -1019 2064
rect -1159 2000 -1019 2047
rect -961 2047 -929 2064
rect -853 2064 -837 2081
rect -747 2081 -639 2097
rect -747 2064 -731 2081
rect -853 2047 -821 2064
rect -961 2000 -821 2047
rect -763 2047 -731 2064
rect -655 2064 -639 2081
rect -549 2081 -441 2097
rect -549 2064 -533 2081
rect -655 2047 -623 2064
rect -763 2000 -623 2047
rect -565 2047 -533 2064
rect -457 2064 -441 2081
rect -351 2081 -243 2097
rect -351 2064 -335 2081
rect -457 2047 -425 2064
rect -565 2000 -425 2047
rect -367 2047 -335 2064
rect -259 2064 -243 2081
rect -153 2081 -45 2097
rect -153 2064 -137 2081
rect -259 2047 -227 2064
rect -367 2000 -227 2047
rect -169 2047 -137 2064
rect -61 2064 -45 2081
rect 45 2081 153 2097
rect 45 2064 61 2081
rect -61 2047 -29 2064
rect -169 2000 -29 2047
rect 29 2047 61 2064
rect 137 2064 153 2081
rect 243 2081 351 2097
rect 243 2064 259 2081
rect 137 2047 169 2064
rect 29 2000 169 2047
rect 227 2047 259 2064
rect 335 2064 351 2081
rect 441 2081 549 2097
rect 441 2064 457 2081
rect 335 2047 367 2064
rect 227 2000 367 2047
rect 425 2047 457 2064
rect 533 2064 549 2081
rect 639 2081 747 2097
rect 639 2064 655 2081
rect 533 2047 565 2064
rect 425 2000 565 2047
rect 623 2047 655 2064
rect 731 2064 747 2081
rect 837 2081 945 2097
rect 837 2064 853 2081
rect 731 2047 763 2064
rect 623 2000 763 2047
rect 821 2047 853 2064
rect 929 2064 945 2081
rect 1035 2081 1143 2097
rect 1035 2064 1051 2081
rect 929 2047 961 2064
rect 821 2000 961 2047
rect 1019 2047 1051 2064
rect 1127 2064 1143 2081
rect 1233 2081 1341 2097
rect 1233 2064 1249 2081
rect 1127 2047 1159 2064
rect 1019 2000 1159 2047
rect 1217 2047 1249 2064
rect 1325 2064 1341 2081
rect 1431 2081 1539 2097
rect 1431 2064 1447 2081
rect 1325 2047 1357 2064
rect 1217 2000 1357 2047
rect 1415 2047 1447 2064
rect 1523 2064 1539 2081
rect 1629 2081 1737 2097
rect 1629 2064 1645 2081
rect 1523 2047 1555 2064
rect 1415 2000 1555 2047
rect 1613 2047 1645 2064
rect 1721 2064 1737 2081
rect 1827 2081 1935 2097
rect 1827 2064 1843 2081
rect 1721 2047 1753 2064
rect 1613 2000 1753 2047
rect 1811 2047 1843 2064
rect 1919 2064 1935 2081
rect 2025 2081 2133 2097
rect 2025 2064 2041 2081
rect 1919 2047 1951 2064
rect 1811 2000 1951 2047
rect 2009 2047 2041 2064
rect 2117 2064 2133 2081
rect 2223 2081 2331 2097
rect 2223 2064 2239 2081
rect 2117 2047 2149 2064
rect 2009 2000 2149 2047
rect 2207 2047 2239 2064
rect 2315 2064 2331 2081
rect 2421 2081 2529 2097
rect 2421 2064 2437 2081
rect 2315 2047 2347 2064
rect 2207 2000 2347 2047
rect 2405 2047 2437 2064
rect 2513 2064 2529 2081
rect 2619 2081 2727 2097
rect 2619 2064 2635 2081
rect 2513 2047 2545 2064
rect 2405 2000 2545 2047
rect 2603 2047 2635 2064
rect 2711 2064 2727 2081
rect 2817 2081 2925 2097
rect 2817 2064 2833 2081
rect 2711 2047 2743 2064
rect 2603 2000 2743 2047
rect 2801 2047 2833 2064
rect 2909 2064 2925 2081
rect 3015 2081 3123 2097
rect 3015 2064 3031 2081
rect 2909 2047 2941 2064
rect 2801 2000 2941 2047
rect 2999 2047 3031 2064
rect 3107 2064 3123 2081
rect 3107 2047 3139 2064
rect 2999 2000 3139 2047
rect -3139 -2047 -2999 -2000
rect -3139 -2064 -3107 -2047
rect -3123 -2081 -3107 -2064
rect -3031 -2064 -2999 -2047
rect -2941 -2047 -2801 -2000
rect -2941 -2064 -2909 -2047
rect -3031 -2081 -3015 -2064
rect -3123 -2097 -3015 -2081
rect -2925 -2081 -2909 -2064
rect -2833 -2064 -2801 -2047
rect -2743 -2047 -2603 -2000
rect -2743 -2064 -2711 -2047
rect -2833 -2081 -2817 -2064
rect -2925 -2097 -2817 -2081
rect -2727 -2081 -2711 -2064
rect -2635 -2064 -2603 -2047
rect -2545 -2047 -2405 -2000
rect -2545 -2064 -2513 -2047
rect -2635 -2081 -2619 -2064
rect -2727 -2097 -2619 -2081
rect -2529 -2081 -2513 -2064
rect -2437 -2064 -2405 -2047
rect -2347 -2047 -2207 -2000
rect -2347 -2064 -2315 -2047
rect -2437 -2081 -2421 -2064
rect -2529 -2097 -2421 -2081
rect -2331 -2081 -2315 -2064
rect -2239 -2064 -2207 -2047
rect -2149 -2047 -2009 -2000
rect -2149 -2064 -2117 -2047
rect -2239 -2081 -2223 -2064
rect -2331 -2097 -2223 -2081
rect -2133 -2081 -2117 -2064
rect -2041 -2064 -2009 -2047
rect -1951 -2047 -1811 -2000
rect -1951 -2064 -1919 -2047
rect -2041 -2081 -2025 -2064
rect -2133 -2097 -2025 -2081
rect -1935 -2081 -1919 -2064
rect -1843 -2064 -1811 -2047
rect -1753 -2047 -1613 -2000
rect -1753 -2064 -1721 -2047
rect -1843 -2081 -1827 -2064
rect -1935 -2097 -1827 -2081
rect -1737 -2081 -1721 -2064
rect -1645 -2064 -1613 -2047
rect -1555 -2047 -1415 -2000
rect -1555 -2064 -1523 -2047
rect -1645 -2081 -1629 -2064
rect -1737 -2097 -1629 -2081
rect -1539 -2081 -1523 -2064
rect -1447 -2064 -1415 -2047
rect -1357 -2047 -1217 -2000
rect -1357 -2064 -1325 -2047
rect -1447 -2081 -1431 -2064
rect -1539 -2097 -1431 -2081
rect -1341 -2081 -1325 -2064
rect -1249 -2064 -1217 -2047
rect -1159 -2047 -1019 -2000
rect -1159 -2064 -1127 -2047
rect -1249 -2081 -1233 -2064
rect -1341 -2097 -1233 -2081
rect -1143 -2081 -1127 -2064
rect -1051 -2064 -1019 -2047
rect -961 -2047 -821 -2000
rect -961 -2064 -929 -2047
rect -1051 -2081 -1035 -2064
rect -1143 -2097 -1035 -2081
rect -945 -2081 -929 -2064
rect -853 -2064 -821 -2047
rect -763 -2047 -623 -2000
rect -763 -2064 -731 -2047
rect -853 -2081 -837 -2064
rect -945 -2097 -837 -2081
rect -747 -2081 -731 -2064
rect -655 -2064 -623 -2047
rect -565 -2047 -425 -2000
rect -565 -2064 -533 -2047
rect -655 -2081 -639 -2064
rect -747 -2097 -639 -2081
rect -549 -2081 -533 -2064
rect -457 -2064 -425 -2047
rect -367 -2047 -227 -2000
rect -367 -2064 -335 -2047
rect -457 -2081 -441 -2064
rect -549 -2097 -441 -2081
rect -351 -2081 -335 -2064
rect -259 -2064 -227 -2047
rect -169 -2047 -29 -2000
rect -169 -2064 -137 -2047
rect -259 -2081 -243 -2064
rect -351 -2097 -243 -2081
rect -153 -2081 -137 -2064
rect -61 -2064 -29 -2047
rect 29 -2047 169 -2000
rect 29 -2064 61 -2047
rect -61 -2081 -45 -2064
rect -153 -2097 -45 -2081
rect 45 -2081 61 -2064
rect 137 -2064 169 -2047
rect 227 -2047 367 -2000
rect 227 -2064 259 -2047
rect 137 -2081 153 -2064
rect 45 -2097 153 -2081
rect 243 -2081 259 -2064
rect 335 -2064 367 -2047
rect 425 -2047 565 -2000
rect 425 -2064 457 -2047
rect 335 -2081 351 -2064
rect 243 -2097 351 -2081
rect 441 -2081 457 -2064
rect 533 -2064 565 -2047
rect 623 -2047 763 -2000
rect 623 -2064 655 -2047
rect 533 -2081 549 -2064
rect 441 -2097 549 -2081
rect 639 -2081 655 -2064
rect 731 -2064 763 -2047
rect 821 -2047 961 -2000
rect 821 -2064 853 -2047
rect 731 -2081 747 -2064
rect 639 -2097 747 -2081
rect 837 -2081 853 -2064
rect 929 -2064 961 -2047
rect 1019 -2047 1159 -2000
rect 1019 -2064 1051 -2047
rect 929 -2081 945 -2064
rect 837 -2097 945 -2081
rect 1035 -2081 1051 -2064
rect 1127 -2064 1159 -2047
rect 1217 -2047 1357 -2000
rect 1217 -2064 1249 -2047
rect 1127 -2081 1143 -2064
rect 1035 -2097 1143 -2081
rect 1233 -2081 1249 -2064
rect 1325 -2064 1357 -2047
rect 1415 -2047 1555 -2000
rect 1415 -2064 1447 -2047
rect 1325 -2081 1341 -2064
rect 1233 -2097 1341 -2081
rect 1431 -2081 1447 -2064
rect 1523 -2064 1555 -2047
rect 1613 -2047 1753 -2000
rect 1613 -2064 1645 -2047
rect 1523 -2081 1539 -2064
rect 1431 -2097 1539 -2081
rect 1629 -2081 1645 -2064
rect 1721 -2064 1753 -2047
rect 1811 -2047 1951 -2000
rect 1811 -2064 1843 -2047
rect 1721 -2081 1737 -2064
rect 1629 -2097 1737 -2081
rect 1827 -2081 1843 -2064
rect 1919 -2064 1951 -2047
rect 2009 -2047 2149 -2000
rect 2009 -2064 2041 -2047
rect 1919 -2081 1935 -2064
rect 1827 -2097 1935 -2081
rect 2025 -2081 2041 -2064
rect 2117 -2064 2149 -2047
rect 2207 -2047 2347 -2000
rect 2207 -2064 2239 -2047
rect 2117 -2081 2133 -2064
rect 2025 -2097 2133 -2081
rect 2223 -2081 2239 -2064
rect 2315 -2064 2347 -2047
rect 2405 -2047 2545 -2000
rect 2405 -2064 2437 -2047
rect 2315 -2081 2331 -2064
rect 2223 -2097 2331 -2081
rect 2421 -2081 2437 -2064
rect 2513 -2064 2545 -2047
rect 2603 -2047 2743 -2000
rect 2603 -2064 2635 -2047
rect 2513 -2081 2529 -2064
rect 2421 -2097 2529 -2081
rect 2619 -2081 2635 -2064
rect 2711 -2064 2743 -2047
rect 2801 -2047 2941 -2000
rect 2801 -2064 2833 -2047
rect 2711 -2081 2727 -2064
rect 2619 -2097 2727 -2081
rect 2817 -2081 2833 -2064
rect 2909 -2064 2941 -2047
rect 2999 -2047 3139 -2000
rect 2999 -2064 3031 -2047
rect 2909 -2081 2925 -2064
rect 2817 -2097 2925 -2081
rect 3015 -2081 3031 -2064
rect 3107 -2064 3139 -2047
rect 3107 -2081 3123 -2064
rect 3015 -2097 3123 -2081
<< polycont >>
rect -3107 2047 -3031 2081
rect -2909 2047 -2833 2081
rect -2711 2047 -2635 2081
rect -2513 2047 -2437 2081
rect -2315 2047 -2239 2081
rect -2117 2047 -2041 2081
rect -1919 2047 -1843 2081
rect -1721 2047 -1645 2081
rect -1523 2047 -1447 2081
rect -1325 2047 -1249 2081
rect -1127 2047 -1051 2081
rect -929 2047 -853 2081
rect -731 2047 -655 2081
rect -533 2047 -457 2081
rect -335 2047 -259 2081
rect -137 2047 -61 2081
rect 61 2047 137 2081
rect 259 2047 335 2081
rect 457 2047 533 2081
rect 655 2047 731 2081
rect 853 2047 929 2081
rect 1051 2047 1127 2081
rect 1249 2047 1325 2081
rect 1447 2047 1523 2081
rect 1645 2047 1721 2081
rect 1843 2047 1919 2081
rect 2041 2047 2117 2081
rect 2239 2047 2315 2081
rect 2437 2047 2513 2081
rect 2635 2047 2711 2081
rect 2833 2047 2909 2081
rect 3031 2047 3107 2081
rect -3107 -2081 -3031 -2047
rect -2909 -2081 -2833 -2047
rect -2711 -2081 -2635 -2047
rect -2513 -2081 -2437 -2047
rect -2315 -2081 -2239 -2047
rect -2117 -2081 -2041 -2047
rect -1919 -2081 -1843 -2047
rect -1721 -2081 -1645 -2047
rect -1523 -2081 -1447 -2047
rect -1325 -2081 -1249 -2047
rect -1127 -2081 -1051 -2047
rect -929 -2081 -853 -2047
rect -731 -2081 -655 -2047
rect -533 -2081 -457 -2047
rect -335 -2081 -259 -2047
rect -137 -2081 -61 -2047
rect 61 -2081 137 -2047
rect 259 -2081 335 -2047
rect 457 -2081 533 -2047
rect 655 -2081 731 -2047
rect 853 -2081 929 -2047
rect 1051 -2081 1127 -2047
rect 1249 -2081 1325 -2047
rect 1447 -2081 1523 -2047
rect 1645 -2081 1721 -2047
rect 1843 -2081 1919 -2047
rect 2041 -2081 2117 -2047
rect 2239 -2081 2315 -2047
rect 2437 -2081 2513 -2047
rect 2635 -2081 2711 -2047
rect 2833 -2081 2909 -2047
rect 3031 -2081 3107 -2047
<< locali >>
rect -3299 2149 -2285 2183
rect 2285 2149 3299 2183
rect -3299 1504 -3265 2149
rect 3265 1504 3299 2149
rect -3185 1392 -3151 1408
rect -3185 -1408 -3151 -1392
rect -2987 1392 -2953 1408
rect -2987 -1408 -2953 -1392
rect -2789 1392 -2755 1408
rect -2789 -1408 -2755 -1392
rect -2591 1392 -2557 1408
rect -2591 -1408 -2557 -1392
rect -2393 1392 -2359 1408
rect -2393 -1408 -2359 -1392
rect -2195 1392 -2161 1408
rect -2195 -1408 -2161 -1392
rect -1997 1392 -1963 1408
rect -1997 -1408 -1963 -1392
rect -1799 1392 -1765 1408
rect -1799 -1408 -1765 -1392
rect -1601 1392 -1567 1408
rect -1601 -1408 -1567 -1392
rect -1403 1392 -1369 1408
rect -1403 -1408 -1369 -1392
rect -1205 1392 -1171 1408
rect -1205 -1408 -1171 -1392
rect -1007 1392 -973 1408
rect -1007 -1408 -973 -1392
rect -809 1392 -775 1408
rect -809 -1408 -775 -1392
rect -611 1392 -577 1408
rect -611 -1408 -577 -1392
rect -413 1392 -379 1408
rect -413 -1408 -379 -1392
rect -215 1392 -181 1408
rect -215 -1408 -181 -1392
rect -17 1392 17 1408
rect -17 -1408 17 -1392
rect 181 1392 215 1408
rect 181 -1408 215 -1392
rect 379 1392 413 1408
rect 379 -1408 413 -1392
rect 577 1392 611 1408
rect 577 -1408 611 -1392
rect 775 1392 809 1408
rect 775 -1408 809 -1392
rect 973 1392 1007 1408
rect 973 -1408 1007 -1392
rect 1171 1392 1205 1408
rect 1171 -1408 1205 -1392
rect 1369 1392 1403 1408
rect 1369 -1408 1403 -1392
rect 1567 1392 1601 1408
rect 1567 -1408 1601 -1392
rect 1765 1392 1799 1408
rect 1765 -1408 1799 -1392
rect 1963 1392 1997 1408
rect 1963 -1408 1997 -1392
rect 2161 1392 2195 1408
rect 2161 -1408 2195 -1392
rect 2359 1392 2393 1408
rect 2359 -1408 2393 -1392
rect 2557 1392 2591 1408
rect 2557 -1408 2591 -1392
rect 2755 1392 2789 1408
rect 2755 -1408 2789 -1392
rect 2953 1392 2987 1408
rect 2953 -1408 2987 -1392
rect 3151 1392 3185 1408
rect 3151 -1408 3185 -1392
rect -3299 -2149 -3265 -1504
rect 3265 -2149 3299 -1504
rect -3299 -2183 -2285 -2149
rect 2285 -2183 3299 -2149
<< viali >>
rect -2285 2149 -2242 2183
rect -2242 2149 2242 2183
rect 2242 2149 2285 2183
rect -3123 2047 -3107 2081
rect -3107 2047 -3031 2081
rect -3031 2047 -3015 2081
rect -2925 2047 -2909 2081
rect -2909 2047 -2833 2081
rect -2833 2047 -2817 2081
rect -2727 2047 -2711 2081
rect -2711 2047 -2635 2081
rect -2635 2047 -2619 2081
rect -2529 2047 -2513 2081
rect -2513 2047 -2437 2081
rect -2437 2047 -2421 2081
rect -2331 2047 -2315 2081
rect -2315 2047 -2239 2081
rect -2239 2047 -2223 2081
rect -2133 2047 -2117 2081
rect -2117 2047 -2041 2081
rect -2041 2047 -2025 2081
rect -1935 2047 -1919 2081
rect -1919 2047 -1843 2081
rect -1843 2047 -1827 2081
rect -1737 2047 -1721 2081
rect -1721 2047 -1645 2081
rect -1645 2047 -1629 2081
rect -1539 2047 -1523 2081
rect -1523 2047 -1447 2081
rect -1447 2047 -1431 2081
rect -1341 2047 -1325 2081
rect -1325 2047 -1249 2081
rect -1249 2047 -1233 2081
rect -1143 2047 -1127 2081
rect -1127 2047 -1051 2081
rect -1051 2047 -1035 2081
rect -945 2047 -929 2081
rect -929 2047 -853 2081
rect -853 2047 -837 2081
rect -747 2047 -731 2081
rect -731 2047 -655 2081
rect -655 2047 -639 2081
rect -549 2047 -533 2081
rect -533 2047 -457 2081
rect -457 2047 -441 2081
rect -351 2047 -335 2081
rect -335 2047 -259 2081
rect -259 2047 -243 2081
rect -153 2047 -137 2081
rect -137 2047 -61 2081
rect -61 2047 -45 2081
rect 45 2047 61 2081
rect 61 2047 137 2081
rect 137 2047 153 2081
rect 243 2047 259 2081
rect 259 2047 335 2081
rect 335 2047 351 2081
rect 441 2047 457 2081
rect 457 2047 533 2081
rect 533 2047 549 2081
rect 639 2047 655 2081
rect 655 2047 731 2081
rect 731 2047 747 2081
rect 837 2047 853 2081
rect 853 2047 929 2081
rect 929 2047 945 2081
rect 1035 2047 1051 2081
rect 1051 2047 1127 2081
rect 1127 2047 1143 2081
rect 1233 2047 1249 2081
rect 1249 2047 1325 2081
rect 1325 2047 1341 2081
rect 1431 2047 1447 2081
rect 1447 2047 1523 2081
rect 1523 2047 1539 2081
rect 1629 2047 1645 2081
rect 1645 2047 1721 2081
rect 1721 2047 1737 2081
rect 1827 2047 1843 2081
rect 1843 2047 1919 2081
rect 1919 2047 1935 2081
rect 2025 2047 2041 2081
rect 2041 2047 2117 2081
rect 2117 2047 2133 2081
rect 2223 2047 2239 2081
rect 2239 2047 2315 2081
rect 2315 2047 2331 2081
rect 2421 2047 2437 2081
rect 2437 2047 2513 2081
rect 2513 2047 2529 2081
rect 2619 2047 2635 2081
rect 2635 2047 2711 2081
rect 2711 2047 2727 2081
rect 2817 2047 2833 2081
rect 2833 2047 2909 2081
rect 2909 2047 2925 2081
rect 3015 2047 3031 2081
rect 3031 2047 3107 2081
rect 3107 2047 3123 2081
rect -3299 1461 -3265 1504
rect -3299 -1461 -3265 1461
rect 3265 1461 3299 1504
rect -3185 -1392 -3151 1392
rect -2987 -1392 -2953 1392
rect -2789 -1392 -2755 1392
rect -2591 -1392 -2557 1392
rect -2393 -1392 -2359 1392
rect -2195 -1392 -2161 1392
rect -1997 -1392 -1963 1392
rect -1799 -1392 -1765 1392
rect -1601 -1392 -1567 1392
rect -1403 -1392 -1369 1392
rect -1205 -1392 -1171 1392
rect -1007 -1392 -973 1392
rect -809 -1392 -775 1392
rect -611 -1392 -577 1392
rect -413 -1392 -379 1392
rect -215 -1392 -181 1392
rect -17 -1392 17 1392
rect 181 -1392 215 1392
rect 379 -1392 413 1392
rect 577 -1392 611 1392
rect 775 -1392 809 1392
rect 973 -1392 1007 1392
rect 1171 -1392 1205 1392
rect 1369 -1392 1403 1392
rect 1567 -1392 1601 1392
rect 1765 -1392 1799 1392
rect 1963 -1392 1997 1392
rect 2161 -1392 2195 1392
rect 2359 -1392 2393 1392
rect 2557 -1392 2591 1392
rect 2755 -1392 2789 1392
rect 2953 -1392 2987 1392
rect 3151 -1392 3185 1392
rect -3299 -1504 -3265 -1461
rect 3265 -1461 3299 1461
rect 3265 -1504 3299 -1461
rect -3123 -2081 -3107 -2047
rect -3107 -2081 -3031 -2047
rect -3031 -2081 -3015 -2047
rect -2925 -2081 -2909 -2047
rect -2909 -2081 -2833 -2047
rect -2833 -2081 -2817 -2047
rect -2727 -2081 -2711 -2047
rect -2711 -2081 -2635 -2047
rect -2635 -2081 -2619 -2047
rect -2529 -2081 -2513 -2047
rect -2513 -2081 -2437 -2047
rect -2437 -2081 -2421 -2047
rect -2331 -2081 -2315 -2047
rect -2315 -2081 -2239 -2047
rect -2239 -2081 -2223 -2047
rect -2133 -2081 -2117 -2047
rect -2117 -2081 -2041 -2047
rect -2041 -2081 -2025 -2047
rect -1935 -2081 -1919 -2047
rect -1919 -2081 -1843 -2047
rect -1843 -2081 -1827 -2047
rect -1737 -2081 -1721 -2047
rect -1721 -2081 -1645 -2047
rect -1645 -2081 -1629 -2047
rect -1539 -2081 -1523 -2047
rect -1523 -2081 -1447 -2047
rect -1447 -2081 -1431 -2047
rect -1341 -2081 -1325 -2047
rect -1325 -2081 -1249 -2047
rect -1249 -2081 -1233 -2047
rect -1143 -2081 -1127 -2047
rect -1127 -2081 -1051 -2047
rect -1051 -2081 -1035 -2047
rect -945 -2081 -929 -2047
rect -929 -2081 -853 -2047
rect -853 -2081 -837 -2047
rect -747 -2081 -731 -2047
rect -731 -2081 -655 -2047
rect -655 -2081 -639 -2047
rect -549 -2081 -533 -2047
rect -533 -2081 -457 -2047
rect -457 -2081 -441 -2047
rect -351 -2081 -335 -2047
rect -335 -2081 -259 -2047
rect -259 -2081 -243 -2047
rect -153 -2081 -137 -2047
rect -137 -2081 -61 -2047
rect -61 -2081 -45 -2047
rect 45 -2081 61 -2047
rect 61 -2081 137 -2047
rect 137 -2081 153 -2047
rect 243 -2081 259 -2047
rect 259 -2081 335 -2047
rect 335 -2081 351 -2047
rect 441 -2081 457 -2047
rect 457 -2081 533 -2047
rect 533 -2081 549 -2047
rect 639 -2081 655 -2047
rect 655 -2081 731 -2047
rect 731 -2081 747 -2047
rect 837 -2081 853 -2047
rect 853 -2081 929 -2047
rect 929 -2081 945 -2047
rect 1035 -2081 1051 -2047
rect 1051 -2081 1127 -2047
rect 1127 -2081 1143 -2047
rect 1233 -2081 1249 -2047
rect 1249 -2081 1325 -2047
rect 1325 -2081 1341 -2047
rect 1431 -2081 1447 -2047
rect 1447 -2081 1523 -2047
rect 1523 -2081 1539 -2047
rect 1629 -2081 1645 -2047
rect 1645 -2081 1721 -2047
rect 1721 -2081 1737 -2047
rect 1827 -2081 1843 -2047
rect 1843 -2081 1919 -2047
rect 1919 -2081 1935 -2047
rect 2025 -2081 2041 -2047
rect 2041 -2081 2117 -2047
rect 2117 -2081 2133 -2047
rect 2223 -2081 2239 -2047
rect 2239 -2081 2315 -2047
rect 2315 -2081 2331 -2047
rect 2421 -2081 2437 -2047
rect 2437 -2081 2513 -2047
rect 2513 -2081 2529 -2047
rect 2619 -2081 2635 -2047
rect 2635 -2081 2711 -2047
rect 2711 -2081 2727 -2047
rect 2817 -2081 2833 -2047
rect 2833 -2081 2909 -2047
rect 2909 -2081 2925 -2047
rect 3015 -2081 3031 -2047
rect 3031 -2081 3107 -2047
rect 3107 -2081 3123 -2047
rect -2285 -2183 -2242 -2149
rect -2242 -2183 2242 -2149
rect 2242 -2183 2285 -2149
<< metal1 >>
rect -2297 2183 2297 2189
rect -2297 2149 -2285 2183
rect 2285 2149 2297 2183
rect -2297 2143 2297 2149
rect -3135 2081 -3003 2087
rect -3135 2047 -3123 2081
rect -3015 2047 -3003 2081
rect -3135 2041 -3003 2047
rect -2937 2081 -2805 2087
rect -2937 2047 -2925 2081
rect -2817 2047 -2805 2081
rect -2937 2041 -2805 2047
rect -2739 2081 -2607 2087
rect -2739 2047 -2727 2081
rect -2619 2047 -2607 2081
rect -2739 2041 -2607 2047
rect -2541 2081 -2409 2087
rect -2541 2047 -2529 2081
rect -2421 2047 -2409 2081
rect -2541 2041 -2409 2047
rect -2343 2081 -2211 2087
rect -2343 2047 -2331 2081
rect -2223 2047 -2211 2081
rect -2343 2041 -2211 2047
rect -2145 2081 -2013 2087
rect -2145 2047 -2133 2081
rect -2025 2047 -2013 2081
rect -2145 2041 -2013 2047
rect -1947 2081 -1815 2087
rect -1947 2047 -1935 2081
rect -1827 2047 -1815 2081
rect -1947 2041 -1815 2047
rect -1749 2081 -1617 2087
rect -1749 2047 -1737 2081
rect -1629 2047 -1617 2081
rect -1749 2041 -1617 2047
rect -1551 2081 -1419 2087
rect -1551 2047 -1539 2081
rect -1431 2047 -1419 2081
rect -1551 2041 -1419 2047
rect -1353 2081 -1221 2087
rect -1353 2047 -1341 2081
rect -1233 2047 -1221 2081
rect -1353 2041 -1221 2047
rect -1155 2081 -1023 2087
rect -1155 2047 -1143 2081
rect -1035 2047 -1023 2081
rect -1155 2041 -1023 2047
rect -957 2081 -825 2087
rect -957 2047 -945 2081
rect -837 2047 -825 2081
rect -957 2041 -825 2047
rect -759 2081 -627 2087
rect -759 2047 -747 2081
rect -639 2047 -627 2081
rect -759 2041 -627 2047
rect -561 2081 -429 2087
rect -561 2047 -549 2081
rect -441 2047 -429 2081
rect -561 2041 -429 2047
rect -363 2081 -231 2087
rect -363 2047 -351 2081
rect -243 2047 -231 2081
rect -363 2041 -231 2047
rect -165 2081 -33 2087
rect -165 2047 -153 2081
rect -45 2047 -33 2081
rect -165 2041 -33 2047
rect 33 2081 165 2087
rect 33 2047 45 2081
rect 153 2047 165 2081
rect 33 2041 165 2047
rect 231 2081 363 2087
rect 231 2047 243 2081
rect 351 2047 363 2081
rect 231 2041 363 2047
rect 429 2081 561 2087
rect 429 2047 441 2081
rect 549 2047 561 2081
rect 429 2041 561 2047
rect 627 2081 759 2087
rect 627 2047 639 2081
rect 747 2047 759 2081
rect 627 2041 759 2047
rect 825 2081 957 2087
rect 825 2047 837 2081
rect 945 2047 957 2081
rect 825 2041 957 2047
rect 1023 2081 1155 2087
rect 1023 2047 1035 2081
rect 1143 2047 1155 2081
rect 1023 2041 1155 2047
rect 1221 2081 1353 2087
rect 1221 2047 1233 2081
rect 1341 2047 1353 2081
rect 1221 2041 1353 2047
rect 1419 2081 1551 2087
rect 1419 2047 1431 2081
rect 1539 2047 1551 2081
rect 1419 2041 1551 2047
rect 1617 2081 1749 2087
rect 1617 2047 1629 2081
rect 1737 2047 1749 2081
rect 1617 2041 1749 2047
rect 1815 2081 1947 2087
rect 1815 2047 1827 2081
rect 1935 2047 1947 2081
rect 1815 2041 1947 2047
rect 2013 2081 2145 2087
rect 2013 2047 2025 2081
rect 2133 2047 2145 2081
rect 2013 2041 2145 2047
rect 2211 2081 2343 2087
rect 2211 2047 2223 2081
rect 2331 2047 2343 2081
rect 2211 2041 2343 2047
rect 2409 2081 2541 2087
rect 2409 2047 2421 2081
rect 2529 2047 2541 2081
rect 2409 2041 2541 2047
rect 2607 2081 2739 2087
rect 2607 2047 2619 2081
rect 2727 2047 2739 2081
rect 2607 2041 2739 2047
rect 2805 2081 2937 2087
rect 2805 2047 2817 2081
rect 2925 2047 2937 2081
rect 2805 2041 2937 2047
rect 3003 2081 3135 2087
rect 3003 2047 3015 2081
rect 3123 2047 3135 2081
rect 3003 2041 3135 2047
rect -3305 1504 -3259 1516
rect -3305 -1504 -3299 1504
rect -3265 -1504 -3259 1504
rect 3259 1504 3305 1516
rect -3191 1392 -3145 1404
rect -3191 -1392 -3185 1392
rect -3151 -1392 -3145 1392
rect -3191 -1404 -3145 -1392
rect -2993 1392 -2947 1404
rect -2993 -1392 -2987 1392
rect -2953 -1392 -2947 1392
rect -2993 -1404 -2947 -1392
rect -2795 1392 -2749 1404
rect -2795 -1392 -2789 1392
rect -2755 -1392 -2749 1392
rect -2795 -1404 -2749 -1392
rect -2597 1392 -2551 1404
rect -2597 -1392 -2591 1392
rect -2557 -1392 -2551 1392
rect -2597 -1404 -2551 -1392
rect -2399 1392 -2353 1404
rect -2399 -1392 -2393 1392
rect -2359 -1392 -2353 1392
rect -2399 -1404 -2353 -1392
rect -2201 1392 -2155 1404
rect -2201 -1392 -2195 1392
rect -2161 -1392 -2155 1392
rect -2201 -1404 -2155 -1392
rect -2003 1392 -1957 1404
rect -2003 -1392 -1997 1392
rect -1963 -1392 -1957 1392
rect -2003 -1404 -1957 -1392
rect -1805 1392 -1759 1404
rect -1805 -1392 -1799 1392
rect -1765 -1392 -1759 1392
rect -1805 -1404 -1759 -1392
rect -1607 1392 -1561 1404
rect -1607 -1392 -1601 1392
rect -1567 -1392 -1561 1392
rect -1607 -1404 -1561 -1392
rect -1409 1392 -1363 1404
rect -1409 -1392 -1403 1392
rect -1369 -1392 -1363 1392
rect -1409 -1404 -1363 -1392
rect -1211 1392 -1165 1404
rect -1211 -1392 -1205 1392
rect -1171 -1392 -1165 1392
rect -1211 -1404 -1165 -1392
rect -1013 1392 -967 1404
rect -1013 -1392 -1007 1392
rect -973 -1392 -967 1392
rect -1013 -1404 -967 -1392
rect -815 1392 -769 1404
rect -815 -1392 -809 1392
rect -775 -1392 -769 1392
rect -815 -1404 -769 -1392
rect -617 1392 -571 1404
rect -617 -1392 -611 1392
rect -577 -1392 -571 1392
rect -617 -1404 -571 -1392
rect -419 1392 -373 1404
rect -419 -1392 -413 1392
rect -379 -1392 -373 1392
rect -419 -1404 -373 -1392
rect -221 1392 -175 1404
rect -221 -1392 -215 1392
rect -181 -1392 -175 1392
rect -221 -1404 -175 -1392
rect -23 1392 23 1404
rect -23 -1392 -17 1392
rect 17 -1392 23 1392
rect -23 -1404 23 -1392
rect 175 1392 221 1404
rect 175 -1392 181 1392
rect 215 -1392 221 1392
rect 175 -1404 221 -1392
rect 373 1392 419 1404
rect 373 -1392 379 1392
rect 413 -1392 419 1392
rect 373 -1404 419 -1392
rect 571 1392 617 1404
rect 571 -1392 577 1392
rect 611 -1392 617 1392
rect 571 -1404 617 -1392
rect 769 1392 815 1404
rect 769 -1392 775 1392
rect 809 -1392 815 1392
rect 769 -1404 815 -1392
rect 967 1392 1013 1404
rect 967 -1392 973 1392
rect 1007 -1392 1013 1392
rect 967 -1404 1013 -1392
rect 1165 1392 1211 1404
rect 1165 -1392 1171 1392
rect 1205 -1392 1211 1392
rect 1165 -1404 1211 -1392
rect 1363 1392 1409 1404
rect 1363 -1392 1369 1392
rect 1403 -1392 1409 1392
rect 1363 -1404 1409 -1392
rect 1561 1392 1607 1404
rect 1561 -1392 1567 1392
rect 1601 -1392 1607 1392
rect 1561 -1404 1607 -1392
rect 1759 1392 1805 1404
rect 1759 -1392 1765 1392
rect 1799 -1392 1805 1392
rect 1759 -1404 1805 -1392
rect 1957 1392 2003 1404
rect 1957 -1392 1963 1392
rect 1997 -1392 2003 1392
rect 1957 -1404 2003 -1392
rect 2155 1392 2201 1404
rect 2155 -1392 2161 1392
rect 2195 -1392 2201 1392
rect 2155 -1404 2201 -1392
rect 2353 1392 2399 1404
rect 2353 -1392 2359 1392
rect 2393 -1392 2399 1392
rect 2353 -1404 2399 -1392
rect 2551 1392 2597 1404
rect 2551 -1392 2557 1392
rect 2591 -1392 2597 1392
rect 2551 -1404 2597 -1392
rect 2749 1392 2795 1404
rect 2749 -1392 2755 1392
rect 2789 -1392 2795 1392
rect 2749 -1404 2795 -1392
rect 2947 1392 2993 1404
rect 2947 -1392 2953 1392
rect 2987 -1392 2993 1392
rect 2947 -1404 2993 -1392
rect 3145 1392 3191 1404
rect 3145 -1392 3151 1392
rect 3185 -1392 3191 1392
rect 3145 -1404 3191 -1392
rect -3305 -1516 -3259 -1504
rect 3259 -1504 3265 1504
rect 3299 -1504 3305 1504
rect 3259 -1516 3305 -1504
rect -3135 -2047 -3003 -2041
rect -3135 -2081 -3123 -2047
rect -3015 -2081 -3003 -2047
rect -3135 -2087 -3003 -2081
rect -2937 -2047 -2805 -2041
rect -2937 -2081 -2925 -2047
rect -2817 -2081 -2805 -2047
rect -2937 -2087 -2805 -2081
rect -2739 -2047 -2607 -2041
rect -2739 -2081 -2727 -2047
rect -2619 -2081 -2607 -2047
rect -2739 -2087 -2607 -2081
rect -2541 -2047 -2409 -2041
rect -2541 -2081 -2529 -2047
rect -2421 -2081 -2409 -2047
rect -2541 -2087 -2409 -2081
rect -2343 -2047 -2211 -2041
rect -2343 -2081 -2331 -2047
rect -2223 -2081 -2211 -2047
rect -2343 -2087 -2211 -2081
rect -2145 -2047 -2013 -2041
rect -2145 -2081 -2133 -2047
rect -2025 -2081 -2013 -2047
rect -2145 -2087 -2013 -2081
rect -1947 -2047 -1815 -2041
rect -1947 -2081 -1935 -2047
rect -1827 -2081 -1815 -2047
rect -1947 -2087 -1815 -2081
rect -1749 -2047 -1617 -2041
rect -1749 -2081 -1737 -2047
rect -1629 -2081 -1617 -2047
rect -1749 -2087 -1617 -2081
rect -1551 -2047 -1419 -2041
rect -1551 -2081 -1539 -2047
rect -1431 -2081 -1419 -2047
rect -1551 -2087 -1419 -2081
rect -1353 -2047 -1221 -2041
rect -1353 -2081 -1341 -2047
rect -1233 -2081 -1221 -2047
rect -1353 -2087 -1221 -2081
rect -1155 -2047 -1023 -2041
rect -1155 -2081 -1143 -2047
rect -1035 -2081 -1023 -2047
rect -1155 -2087 -1023 -2081
rect -957 -2047 -825 -2041
rect -957 -2081 -945 -2047
rect -837 -2081 -825 -2047
rect -957 -2087 -825 -2081
rect -759 -2047 -627 -2041
rect -759 -2081 -747 -2047
rect -639 -2081 -627 -2047
rect -759 -2087 -627 -2081
rect -561 -2047 -429 -2041
rect -561 -2081 -549 -2047
rect -441 -2081 -429 -2047
rect -561 -2087 -429 -2081
rect -363 -2047 -231 -2041
rect -363 -2081 -351 -2047
rect -243 -2081 -231 -2047
rect -363 -2087 -231 -2081
rect -165 -2047 -33 -2041
rect -165 -2081 -153 -2047
rect -45 -2081 -33 -2047
rect -165 -2087 -33 -2081
rect 33 -2047 165 -2041
rect 33 -2081 45 -2047
rect 153 -2081 165 -2047
rect 33 -2087 165 -2081
rect 231 -2047 363 -2041
rect 231 -2081 243 -2047
rect 351 -2081 363 -2047
rect 231 -2087 363 -2081
rect 429 -2047 561 -2041
rect 429 -2081 441 -2047
rect 549 -2081 561 -2047
rect 429 -2087 561 -2081
rect 627 -2047 759 -2041
rect 627 -2081 639 -2047
rect 747 -2081 759 -2047
rect 627 -2087 759 -2081
rect 825 -2047 957 -2041
rect 825 -2081 837 -2047
rect 945 -2081 957 -2047
rect 825 -2087 957 -2081
rect 1023 -2047 1155 -2041
rect 1023 -2081 1035 -2047
rect 1143 -2081 1155 -2047
rect 1023 -2087 1155 -2081
rect 1221 -2047 1353 -2041
rect 1221 -2081 1233 -2047
rect 1341 -2081 1353 -2047
rect 1221 -2087 1353 -2081
rect 1419 -2047 1551 -2041
rect 1419 -2081 1431 -2047
rect 1539 -2081 1551 -2047
rect 1419 -2087 1551 -2081
rect 1617 -2047 1749 -2041
rect 1617 -2081 1629 -2047
rect 1737 -2081 1749 -2047
rect 1617 -2087 1749 -2081
rect 1815 -2047 1947 -2041
rect 1815 -2081 1827 -2047
rect 1935 -2081 1947 -2047
rect 1815 -2087 1947 -2081
rect 2013 -2047 2145 -2041
rect 2013 -2081 2025 -2047
rect 2133 -2081 2145 -2047
rect 2013 -2087 2145 -2081
rect 2211 -2047 2343 -2041
rect 2211 -2081 2223 -2047
rect 2331 -2081 2343 -2047
rect 2211 -2087 2343 -2081
rect 2409 -2047 2541 -2041
rect 2409 -2081 2421 -2047
rect 2529 -2081 2541 -2047
rect 2409 -2087 2541 -2081
rect 2607 -2047 2739 -2041
rect 2607 -2081 2619 -2047
rect 2727 -2081 2739 -2047
rect 2607 -2087 2739 -2081
rect 2805 -2047 2937 -2041
rect 2805 -2081 2817 -2047
rect 2925 -2081 2937 -2047
rect 2805 -2087 2937 -2081
rect 3003 -2047 3135 -2041
rect 3003 -2081 3015 -2047
rect 3123 -2081 3135 -2047
rect 3003 -2087 3135 -2081
rect -2297 -2149 2297 -2143
rect -2297 -2183 -2285 -2149
rect 2285 -2183 2297 -2149
rect -2297 -2189 2297 -2183
<< properties >>
string FIXED_BBOX -3282 -2166 3282 2166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 20.0 l 0.7 m 1 nf 32 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
