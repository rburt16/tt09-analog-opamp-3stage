magic
tech sky130A
magscale 1 2
timestamp 1729530615
<< error_p >>
rect -31 1081 31 1087
rect -31 1047 -19 1081
rect -31 1041 31 1047
rect -31 -1047 31 -1041
rect -31 -1081 -19 -1047
rect -31 -1087 31 -1081
<< nwell >>
rect -231 -1219 231 1219
<< pmoslvt >>
rect -35 -1000 35 1000
<< pdiff >>
rect -93 988 -35 1000
rect -93 -988 -81 988
rect -47 -988 -35 988
rect -93 -1000 -35 -988
rect 35 988 93 1000
rect 35 -988 47 988
rect 81 -988 93 988
rect 35 -1000 93 -988
<< pdiffc >>
rect -81 -988 -47 988
rect 47 -988 81 988
<< nsubdiff >>
rect -195 1149 -99 1183
rect 99 1149 195 1183
rect -195 1087 -161 1149
rect 161 1087 195 1149
rect -195 -1149 -161 -1087
rect 161 -1149 195 -1087
rect -195 -1183 -99 -1149
rect 99 -1183 195 -1149
<< nsubdiffcont >>
rect -99 1149 99 1183
rect -195 -1087 -161 1087
rect 161 -1087 195 1087
rect -99 -1183 99 -1149
<< poly >>
rect -35 1081 35 1097
rect -35 1047 -19 1081
rect 19 1047 35 1081
rect -35 1000 35 1047
rect -35 -1047 35 -1000
rect -35 -1081 -19 -1047
rect 19 -1081 35 -1047
rect -35 -1097 35 -1081
<< polycont >>
rect -19 1047 19 1081
rect -19 -1081 19 -1047
<< locali >>
rect -195 1149 -99 1183
rect 99 1149 195 1183
rect -195 1087 -161 1149
rect 161 1087 195 1149
rect -35 1047 -19 1081
rect 19 1047 35 1081
rect -81 988 -47 1004
rect -81 -1004 -47 -988
rect 47 988 81 1004
rect 47 -1004 81 -988
rect -35 -1081 -19 -1047
rect 19 -1081 35 -1047
rect -195 -1149 -161 -1087
rect 161 -1149 195 -1087
rect -195 -1183 -99 -1149
rect 99 -1183 195 -1149
<< viali >>
rect -19 1047 19 1081
rect -81 -988 -47 988
rect 47 -988 81 988
rect -19 -1081 19 -1047
<< metal1 >>
rect -31 1081 31 1087
rect -31 1047 -19 1081
rect 19 1047 31 1081
rect -31 1041 31 1047
rect -87 988 -41 1000
rect -87 -988 -81 988
rect -47 -988 -41 988
rect -87 -1000 -41 -988
rect 41 988 87 1000
rect 41 -988 47 988
rect 81 -988 87 988
rect 41 -1000 87 -988
rect -31 -1047 31 -1041
rect -31 -1081 -19 -1047
rect 19 -1081 31 -1047
rect -31 -1087 31 -1081
<< properties >>
string FIXED_BBOX -178 -1166 178 1166
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
