* NGSPICE file created from op_amp_3stage.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_M5XJZ4 a_158_n1064# a_358_n1000# a_n358_n1064# a_n158_n1000#
+ a_n416_n1000# a_100_n1000# a_n100_n1064# w_n554_n1219#
X0 a_358_n1000# a_158_n1064# a_100_n1000# w_n554_n1219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X1 a_100_n1000# a_n100_n1064# a_n158_n1000# w_n554_n1219# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X2 a_n158_n1000# a_n358_n1064# a_n416_n1000# w_n554_n1219# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_PP2UM9 a_n458_n1709# a_n400_54# a_n458_109# a_n400_n1764#
+ a_400_n1709# a_400_109# a_n560_n1883#
X0 a_400_109# a_n400_54# a_n458_109# a_n560_n1883# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=4
X1 a_400_n1709# a_n400_n1764# a_n458_n1709# a_n560_n1883# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=4
.ends

.subckt sky130_fd_pr__pfet_01v8_MD8735 a_358_n2118# a_n416_118# a_n158_n2118# a_158_n2182#
+ a_n100_54# a_n358_54# a_358_118# a_158_54# a_n416_n2118# a_n358_n2182# a_n158_118#
+ a_100_n2118# a_n100_n2182# w_n554_n2337# a_100_118#
X0 a_100_118# a_n100_54# a_n158_118# w_n554_n2337# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X1 a_358_n2118# a_158_n2182# a_100_n2118# w_n554_n2337# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X2 a_100_n2118# a_n100_n2182# a_n158_n2118# w_n554_n2337# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X3 a_n158_n2118# a_n358_n2182# a_n416_n2118# w_n554_n2337# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X4 a_358_118# a_158_54# a_100_118# w_n554_n2337# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X5 a_n158_118# a_n358_54# a_n416_118# w_n554_n2337# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_M7ZRRL a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219#
X0 a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_QW8YAA a_n29_n2000# a_29_n2055# a_1629_n2000#
+ a_n1789_n2174# a_n1629_n2055# a_n1687_n2000#
X0 a_1629_n2000# a_29_n2055# a_n29_n2000# a_n1789_n2174# sky130_fd_pr__nfet_01v8_lvt ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=8
X1 a_n29_n2000# a_n1629_n2055# a_n1687_n2000# a_n1789_n2174# sky130_fd_pr__nfet_01v8_lvt ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_WA2NKZ a_n400_n3218# a_n400_n4036# a_n400_n1582#
+ a_n458_n3981# a_n400_54# a_400_927# a_n458_1745# a_n458_2563# a_n458_3381# a_n458_109#
+ a_n400_n2400# a_400_n1527# a_400_n2345# a_400_n3163# a_n400_n764# a_400_n709# a_n458_927#
+ a_n400_2508# a_n400_3326# a_n560_n4155# a_400_n3981# a_n400_1690# a_n458_n1527#
+ a_n458_n709# a_400_109# a_n458_n3163# a_n458_n2345# a_n400_872# a_400_1745# a_400_2563#
+ a_400_3381#
X0 a_400_1745# a_n400_1690# a_n458_1745# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X1 a_400_109# a_n400_54# a_n458_109# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X2 a_400_n1527# a_n400_n1582# a_n458_n1527# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X3 a_400_927# a_n400_872# a_n458_927# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X4 a_400_2563# a_n400_2508# a_n458_2563# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X5 a_400_n2345# a_n400_n2400# a_n458_n2345# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X6 a_400_n709# a_n400_n764# a_n458_n709# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X7 a_400_3381# a_n400_3326# a_n458_3381# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X8 a_400_n3163# a_n400_n3218# a_n458_n3163# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
X9 a_400_n3981# a_n400_n4036# a_n458_n3981# a_n560_n4155# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MXC9RL a_n93_118# a_n35_n2182# a_n93_n2118# a_35_118#
+ a_n35_54# a_35_n2118# w_n231_n2337#
X0 a_35_n2118# a_n35_n2182# a_n93_n2118# w_n231_n2337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1 a_35_118# a_n35_54# a_n93_118# w_n231_n2337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_W9NHZX a_n93_n250# a_n195_n424# a_n35_n305# a_35_n250#
X0 a_35_n250# a_n35_n305# a_n93_n250# a_n195_n424# sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.35
.ends

.subckt sky130_fd_pr__pfet_01v8_L7EPZQ a_100_n836# w_n296_n984# a_n158_n836# a_n100_n862#
X0 a_100_n836# a_n100_n862# a_n158_n836# w_n296_n984# sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_LBMMZQ a_100_n836# w_n296_n984# a_n158_n836# a_n100_n862#
X0 a_100_n836# a_n100_n862# a_n158_n836# w_n296_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_GQTHCS a_800_n78# a_n800_n104# a_n858_n78# w_n996_n226#
X0 a_800_n78# a_n800_n104# a_n858_n78# w_n996_n226# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_N4YVNS a_800_n73# a_n800_n99# a_n858_n73# a_n960_n185#
X0 a_800_n73# a_n800_n99# a_n858_n73# a_n960_n185# sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_QGAK58 a_n158_n831# a_n260_n943# a_100_n831# a_n100_n857#
X0 a_100_n831# a_n100_n857# a_n158_n831# a_n260_n943# sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_BMAEVH a_100_n836# w_n296_n984# a_n158_n836# a_n100_n862#
X0 a_100_n836# a_n100_n862# a_n158_n836# w_n296_n984# sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_92UKLN a_n158_n831# a_n260_n943# a_100_n831# a_n100_n857#
X0 a_100_n831# a_n100_n857# a_n158_n831# a_n260_n943# sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_798YF4 a_n1310_n157# a_1310_n131# a_n1368_n131# a_n1470_n243#
X0 a_1310_n131# a_n1310_n157# a_n1368_n131# a_n1470_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=13.1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_XLZA2Q a_n158_n831# a_n260_n943# a_100_n831# a_n100_n857#
X0 a_100_n831# a_n100_n857# a_n158_n831# a_n260_n943# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_EE6UX6 a_800_n131# a_n800_n157# a_n858_n131# a_n960_n243#
X0 a_800_n131# a_n800_n157# a_n858_n131# a_n960_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_X6KF3T a_n158_n831# a_n260_n943# a_100_n831# a_n100_n857#
X0 a_100_n831# a_n100_n857# a_n158_n831# a_n260_n943# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_LHEPZQ a_100_n836# w_n296_n984# a_n158_n836# a_n100_n862#
X0 a_100_n836# a_n100_n862# a_n158_n836# w_n296_n984# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
.ends

.subckt bias_generator m1_8340_6460# m1_3200_5840# VSUBS
Xsky130_fd_pr__pfet_01v8_L7EPZQ_0 m1_7900_4600# m1_3200_5840# m1_3200_5840# m1_5740_4600#
+ sky130_fd_pr__pfet_01v8_L7EPZQ
XXM12 m1_5740_4600# m1_3200_5840# m1_5260_4600# m1_5740_4600# sky130_fd_pr__pfet_01v8_lvt_LBMMZQ
XXM13 m1_8880_2800# m1_3200_5840# m1_6940_4620# m1_5740_4600# sky130_fd_pr__pfet_01v8_lvt_LBMMZQ
XXM16 m1_9560_5780# m1_3400_4220# m1_3200_5840# m1_3200_5840# sky130_fd_pr__pfet_01v8_GQTHCS
XXM18 VSUBS m1_9560_5780# m1_5740_4600# VSUBS sky130_fd_pr__nfet_01v8_N4YVNS
Xsky130_fd_pr__nfet_01v8_QGAK58_0 m1_9560_5780# VSUBS VSUBS m1_3400_4220# sky130_fd_pr__nfet_01v8_QGAK58
Xsky130_fd_pr__pfet_01v8_lvt_LBMMZQ_0 m1_8340_6460# m1_3200_5840# m1_7900_4600# m1_5740_4600#
+ sky130_fd_pr__pfet_01v8_lvt_LBMMZQ
XXM3 m1_3580_4600# m1_3200_5840# m1_3200_5840# m1_5740_4600# sky130_fd_pr__pfet_01v8_BMAEVH
XXM4 m1_5260_4600# m1_3200_5840# m1_3200_5840# m1_5740_4600# sky130_fd_pr__pfet_01v8_L7EPZQ
XXM6 m1_6940_4620# m1_3200_5840# m1_3200_5840# m1_5740_4600# sky130_fd_pr__pfet_01v8_L7EPZQ
Xsky130_fd_pr__nfet_01v8_92UKLN_1 m1_3400_4220# VSUBS VSUBS m1_3400_4220# sky130_fd_pr__nfet_01v8_92UKLN
Xsky130_fd_pr__nfet_01v8_92UKLN_0 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
XXM7 m1_8880_2800# m1_8880_2800# m1_7680_3620# VSUBS sky130_fd_pr__nfet_01v8_798YF4
Xsky130_fd_pr__nfet_01v8_92UKLN_2 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
XXM9 m1_4380_6140# VSUBS m1_3400_4220# m1_4380_6140# sky130_fd_pr__nfet_01v8_lvt_XLZA2Q
XXM8 m1_3580_2360# m1_8880_2800# m1_7680_3620# VSUBS sky130_fd_pr__nfet_01v8_EE6UX6
Xsky130_fd_pr__nfet_01v8_92UKLN_3 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
Xsky130_fd_pr__nfet_01v8_EE6UX6_1 m1_3580_2360# m1_8880_2800# VSUBS VSUBS sky130_fd_pr__nfet_01v8_EE6UX6
Xsky130_fd_pr__nfet_01v8_EE6UX6_0 m1_3580_2360# m1_8880_2800# VSUBS VSUBS sky130_fd_pr__nfet_01v8_EE6UX6
Xsky130_fd_pr__nfet_01v8_92UKLN_4 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
Xsky130_fd_pr__nfet_01v8_92UKLN_5 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
Xsky130_fd_pr__nfet_01v8_92UKLN_6 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
Xsky130_fd_pr__nfet_01v8_92UKLN_7 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
Xsky130_fd_pr__nfet_01v8_92UKLN_8 m1_3280_4120# VSUBS m1_3580_2360# m1_3400_4220#
+ sky130_fd_pr__nfet_01v8_92UKLN
XXM10 m1_5740_4600# VSUBS m1_3280_4120# m1_4380_6140# sky130_fd_pr__nfet_01v8_lvt_X6KF3T
XXM11 m1_4380_6140# m1_3200_5840# m1_3580_4600# m1_5740_4600# sky130_fd_pr__pfet_01v8_lvt_LHEPZQ
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_545GKL a_367_n2000# a_425_n2064# a_n367_n2064#
+ a_169_n2000# a_n3197_n2000# a_227_n2064# a_n169_n2064# w_n3335_n2219# a_n821_n2000#
+ a_n623_n2000# a_n29_n2000# a_n425_n2000# a_n227_n2000# a_n1951_n2064# a_n2941_n2064#
+ a_2941_n2000# a_n2743_n2064# a_1951_n2000# a_n1753_n2064# a_2743_n2000# a_1753_n2000#
+ a_2801_n2064# a_1811_n2064# a_n1555_n2064# a_n2545_n2064# a_2545_n2000# a_2603_n2064#
+ a_n2347_n2064# a_1555_n2000# a_1613_n2064# a_n1357_n2064# a_n3139_n2064# a_2347_n2000#
+ a_1357_n2000# a_2405_n2064# a_1415_n2064# a_n1159_n2064# a_n2149_n2064# a_3139_n2000#
+ a_2149_n2000# a_1159_n2000# a_2207_n2064# a_1217_n2064# a_n2801_n2000# a_2999_n2064#
+ a_2009_n2064# a_1019_n2064# a_n1811_n2000# a_n1613_n2000# a_n2603_n2000# a_n2405_n2000#
+ a_n1415_n2000# a_n1217_n2000# a_n2207_n2000# a_29_n2064# a_n2009_n2000# a_n2999_n2000#
+ a_961_n2000# a_n1019_n2000# a_n961_n2064# a_763_n2000# a_821_n2064# a_n763_n2064#
+ a_565_n2000# a_623_n2064# a_n565_n2064#
X0 a_1753_n2000# a_1613_n2064# a_1555_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X1 a_n2801_n2000# a_n2941_n2064# a_n2999_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X2 a_367_n2000# a_227_n2064# a_169_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X3 a_n623_n2000# a_n763_n2064# a_n821_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X4 a_n1019_n2000# a_n1159_n2064# a_n1217_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X5 a_1357_n2000# a_1217_n2064# a_1159_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X6 a_n2405_n2000# a_n2545_n2064# a_n2603_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X7 a_2743_n2000# a_2603_n2064# a_2545_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X8 a_n227_n2000# a_n367_n2064# a_n425_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X9 a_961_n2000# a_821_n2064# a_763_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X10 a_n2009_n2000# a_n2149_n2064# a_n2207_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X11 a_2347_n2000# a_2207_n2064# a_2149_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X12 a_n1613_n2000# a_n1753_n2064# a_n1811_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X13 a_1951_n2000# a_1811_n2064# a_1753_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X14 a_565_n2000# a_425_n2064# a_367_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X15 a_n821_n2000# a_n961_n2064# a_n1019_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X16 a_n1217_n2000# a_n1357_n2064# a_n1415_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X17 a_n2999_n2000# a_n3139_n2064# a_n3197_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=5.8 ps=40.58 w=20 l=0.7
X18 a_1555_n2000# a_1415_n2064# a_1357_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X19 a_n2603_n2000# a_n2743_n2064# a_n2801_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X20 a_2941_n2000# a_2801_n2064# a_2743_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X21 a_n425_n2000# a_n565_n2064# a_n623_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X22 a_1159_n2000# a_1019_n2064# a_961_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X23 a_n2207_n2000# a_n2347_n2064# a_n2405_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X24 a_n1811_n2000# a_n1951_n2064# a_n2009_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X25 a_2545_n2000# a_2405_n2064# a_2347_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X26 a_n29_n2000# a_n169_n2064# a_n227_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X27 a_763_n2000# a_623_n2064# a_565_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X28 a_n1415_n2000# a_n1555_n2064# a_n1613_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X29 a_169_n2000# a_29_n2064# a_n29_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X30 a_2149_n2000# a_2009_n2064# a_1951_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.29 as=2.9 ps=20.29 w=20 l=0.7
X31 a_3139_n2000# a_2999_n2064# a_2941_n2000# w_n3335_n2219# sky130_fd_pr__pfet_01v8_lvt ad=5.8 pd=40.58 as=2.9 ps=20.29 w=20 l=0.7
.ends

.subckt sky130_fd_pr__pfet_01v8_M7ZEKL a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219#
X0 a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_C84B7J a_100_n169# a_n260_n343# a_n100_n224# a_n158_n169#
X0 a_100_n169# a_n100_n224# a_n158_n169# a_n260_n343# sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_SHAVFW a_861_n664# a_477_n664# a_803_109# a_n477_109#
+ a_n1059_54# a_803_n609# a_419_n609# a_n349_n609# a_n733_n609# a_n163_n664# a_n733_109#
+ a_163_n609# a_221_54# a_n291_54# a_989_n664# a_221_n664# a_n803_54# a_n93_n609#
+ a_675_109# a_n419_54# a_35_109# a_733_54# a_349_54# a_n675_n664# a_675_n609# a_931_109#
+ a_733_n664# a_n221_109# a_93_54# a_349_n664# a_n605_n609# a_n1117_n609# a_n861_109#
+ a_163_109# a_n35_n664# a_93_n664# a_n931_54# a_35_n609# a_n1117_109# a_n547_54#
+ a_n1219_n783# a_419_109# a_861_54# a_477_54# a_n547_n664# a_n931_n664# a_n1059_n664#
+ a_931_n609# a_1059_109# a_547_n609# a_n861_n609# a_n93_109# a_n477_n609# a_605_n664#
+ a_n349_109# a_989_54# a_n291_n664# a_291_109# a_n605_109# a_n989_109# a_291_n609#
+ a_n35_54# a_n163_54# a_1059_n609# a_n221_n609# a_n989_n609# a_547_109# a_605_54#
+ a_n675_54# a_n419_n664# a_n803_n664#
X0 a_n349_n609# a_n419_n664# a_n477_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X1 a_n861_109# a_n931_54# a_n989_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X2 a_n477_109# a_n547_54# a_n605_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X3 a_n93_109# a_n163_54# a_n221_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X4 a_163_109# a_93_54# a_35_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X5 a_803_n609# a_733_n664# a_675_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X6 a_291_n609# a_221_n664# a_163_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X7 a_803_109# a_733_54# a_675_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X8 a_419_109# a_349_54# a_291_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X9 a_n221_n609# a_n291_n664# a_n349_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X10 a_419_n609# a_349_n664# a_291_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X11 a_n861_n609# a_n931_n664# a_n989_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X12 a_35_n609# a_n35_n664# a_n93_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X13 a_35_109# a_n35_54# a_n93_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X14 a_1059_109# a_989_54# a_931_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.35
X15 a_n477_n609# a_n547_n664# a_n605_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X16 a_n989_n609# a_n1059_n664# a_n1117_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.35
X17 a_931_n609# a_861_n664# a_803_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X18 a_n733_109# a_n803_54# a_n861_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X19 a_n349_109# a_n419_54# a_n477_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X20 a_291_109# a_221_54# a_163_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X21 a_1059_n609# a_989_n664# a_931_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.35
X22 a_675_109# a_605_54# a_547_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X23 a_547_n609# a_477_n664# a_419_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X24 a_n989_109# a_n1059_54# a_n1117_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.35
X25 a_n221_109# a_n291_54# a_n349_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X26 a_163_n609# a_93_n664# a_35_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X27 a_n605_109# a_n675_54# a_n733_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X28 a_675_n609# a_605_n664# a_547_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X29 a_547_109# a_477_54# a_419_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X30 a_931_109# a_861_54# a_803_109# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X31 a_n605_n609# a_n675_n664# a_n733_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X32 a_n93_n609# a_n163_n664# a_n221_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
X33 a_n733_n609# a_n803_n664# a_n861_n609# a_n1219_n783# sky130_fd_pr__nfet_01v8_lvt ad=0.3625 pd=2.79 as=0.3625 ps=2.79 w=2.5 l=0.35
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_QQJVLQ a_163_118# a_419_n2118# a_419_118# a_221_54#
+ a_n291_54# a_n349_n2118# a_349_n2182# a_n733_n2118# a_n675_n2182# a_n93_118# a_n349_118#
+ a_n419_54# a_n291_n2182# a_349_54# a_n35_n2182# a_291_118# a_n605_118# a_93_54#
+ a_93_n2182# a_n419_n2182# a_547_118# a_547_n2118# a_163_n2118# a_n477_118# a_n93_n2118#
+ a_n547_54# a_477_54# a_n477_n2118# a_477_n2182# a_n733_118# a_675_118# w_n871_n2337#
+ a_n605_n2118# a_605_n2182# a_n547_n2182# a_35_118# a_n221_n2118# a_221_n2182# a_n163_n2182#
+ a_n35_54# a_n163_54# a_35_n2118# a_n221_118# a_605_54# a_n675_54# a_675_n2118# a_291_n2118#
X0 a_n221_118# a_n291_54# a_n349_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X1 a_n605_118# a_n675_54# a_n733_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.35
X2 a_291_n2118# a_221_n2182# a_163_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X3 a_419_n2118# a_349_n2182# a_291_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X4 a_547_118# a_477_54# a_419_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X5 a_163_n2118# a_93_n2182# a_35_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X6 a_35_n2118# a_n35_n2182# a_n93_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X7 a_n93_118# a_n163_54# a_n221_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X8 a_163_118# a_93_54# a_35_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X9 a_n477_118# a_n547_54# a_n605_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X10 a_419_118# a_349_54# a_291_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X11 a_n605_n2118# a_n675_n2182# a_n733_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.35
X12 a_n221_n2118# a_n291_n2182# a_n349_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X13 a_35_118# a_n35_54# a_n93_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X14 a_n477_n2118# a_n547_n2182# a_n605_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X15 a_n93_n2118# a_n163_n2182# a_n221_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X16 a_547_n2118# a_477_n2182# a_419_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X17 a_n349_118# a_n419_54# a_n477_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X18 a_291_118# a_221_54# a_163_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
X19 a_675_118# a_605_54# a_547_118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.35
X20 a_675_n2118# a_605_n2182# a_547_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.35
X21 a_n349_n2118# a_n419_n2182# a_n477_n2118# w_n871_n2337# sky130_fd_pr__pfet_01v8_lvt ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_Q53FMB a_n93_n250# a_n195_n424# a_n35_n305# a_35_n250#
X0 a_35_n250# a_n35_n305# a_n93_n250# a_n195_n424# sky130_fd_pr__nfet_01v8_lvt ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.35
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_PD3USF a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219#
X0 a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_SLP2FE a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219#
X0 a_35_n1000# a_n35_n1064# a_n93_n1000# w_n231_n1219# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
.ends

.subckt sky130_fd_pr__pfet_01v8_MV5GT4 a_358_n4354# a_158_n4418# a_358_n2118# a_n416_118#
+ a_n158_n4354# a_n158_n2118# a_158_n2182# a_n100_54# a_n358_54# a_158_2290# a_358_118#
+ a_158_54# a_n358_n4418# a_358_2354# a_n416_n4354# a_n416_n2118# a_n358_n2182# a_n158_118#
+ a_100_2354# a_n358_2290# a_100_n4354# a_100_n2118# a_n158_2354# a_n100_2290# a_n100_n4418#
+ a_n100_n2182# w_n554_n4573# a_100_118# a_n416_2354#
X0 a_100_2354# a_n100_2290# a_n158_2354# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X1 a_100_118# a_n100_54# a_n158_118# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X2 a_358_n4354# a_158_n4418# a_100_n4354# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X3 a_n158_n4354# a_n358_n4418# a_n416_n4354# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X4 a_100_n4354# a_n100_n4418# a_n158_n4354# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X5 a_n158_2354# a_n358_2290# a_n416_2354# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X6 a_358_n2118# a_158_n2182# a_100_n2118# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X7 a_100_n2118# a_n100_n2182# a_n158_n2118# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X8 a_n158_n2118# a_n358_n2182# a_n416_n2118# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X9 a_358_2354# a_158_2290# a_100_2354# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X10 a_358_118# a_158_54# a_100_118# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X11 a_n158_118# a_n358_54# a_n416_118# w_n554_n4573# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_A4BC7Z m3_n2886_n1040# c1_n2846_n1000#
X0 c1_n2846_n1000# m3_n2886_n1040# sky130_fd_pr__cap_mim_m3_1 l=10 w=27
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MF6SRL a_n93_118# a_n35_n4418# a_n35_n2182# a_n93_2354#
+ a_n93_n4354# a_n93_n2118# a_35_2354# a_35_118# a_n35_54# a_35_n4354# a_35_n2118#
+ w_n231_n4573# a_n35_2290#
X0 a_35_n4354# a_n35_n4418# a_n93_n4354# w_n231_n4573# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X1 a_35_2354# a_n35_2290# a_n93_2354# w_n231_n4573# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X2 a_35_n2118# a_n35_n2182# a_n93_n2118# w_n231_n4573# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X3 a_35_118# a_n35_54# a_n93_118# w_n231_n4573# sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_N28DAC a_n560_n474# a_n400_n355# a_400_n300# a_n458_n300#
X0 a_400_n300# a_n400_n355# a_n458_n300# a_n560_n474# sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=4
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_5HBWYY m3_n3186_n2740# c1_n3146_n2700#
X0 c1_n3146_n2700# m3_n3186_n2740# sky130_fd_pr__cap_mim_m3_1 l=27 w=30
.ends

.subckt sky130_fd_pr__pfet_01v8_JHT74A a_n227_n1000# w_n365_n1219# a_29_n1064# a_169_n1000#
+ a_n169_n1064# a_n29_n1000#
X0 a_169_n1000# a_29_n1064# a_n29_n1000# w_n365_n1219# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=0.7
X1 a_n29_n1000# a_n169_n1064# a_n227_n1000# w_n365_n1219# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=0.7
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FWQUH5 a_n458_n800# a_n560_n974# a_n400_n855#
+ a_400_n800#
X0 a_400_n800# a_n400_n855# a_n458_n800# a_n560_n974# sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=4
.ends

.subckt sky130_fd_pr__pfet_01v8_F4HV3A a_n93_n250# a_35_n250# w_n231_n469# a_n35_n314#
X0 a_35_n250# a_n35_n314# a_n93_n250# w_n231_n469# sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=0.35
.ends

.subckt op_amp_3stage
Xsky130_fd_pr__pfet_01v8_M5XJZ4_0 m1_n41520_15180# m1_n41290_29050# m1_n41520_15180#
+ m1_n41290_29050# w_n40780_17110# w_n40780_17110# m1_n41520_15180# w_n40780_17110#
+ sky130_fd_pr__pfet_01v8_M5XJZ4
XXM34 m1_n36990_22880# m1_n37390_15270# m1_n36990_22880# m1_n37390_15270# VSUBS VSUBS
+ VSUBS sky130_fd_pr__nfet_01v8_lvt_PP2UM9
XXM36 m1_n37110_25500# w_n40780_17110# m1_n37110_25500# m1_n41520_15180# m1_n41520_15180#
+ m1_n41520_15180# m1_n37110_25500# m1_n41520_15180# w_n40780_17110# m1_n41520_15180#
+ m1_n37110_25500# w_n40780_17110# m1_n41520_15180# w_n40780_17110# w_n40780_17110#
+ sky130_fd_pr__pfet_01v8_MD8735
XXM35 m1_n40050_29050# m1_n41520_15180# m1_n41290_29050# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_M7ZRRL
XXM14 VSUBS m1_n30380_9040# m4_n35400_n620# VSUBS m1_n30380_9040# m4_n35400_n620#
+ sky130_fd_pr__nfet_01v8_lvt_QW8YAA
XXM25 m1_n41520_15180# m1_n39200_16970# m1_n41520_15180# m1_n39200_16970# w_n40780_17110#
+ w_n40780_17110# m1_n41520_15180# w_n40780_17110# sky130_fd_pr__pfet_01v8_M5XJZ4
XXM24 m1_n33750_9350# m1_n33750_9350# m1_n33750_9350# m1_n33990_17300# m1_n33750_9350#
+ VSUBS m1_n33990_17300# m1_n33990_17300# m1_n33990_17300# m1_n33990_17300# m1_n33750_9350#
+ VSUBS VSUBS VSUBS m1_n33750_9350# VSUBS m1_n33990_17300# m1_n33750_9350# m1_n33750_9350#
+ VSUBS VSUBS m1_n33750_9350# m1_n33990_17300# m1_n33990_17300# VSUBS m1_n33990_17300#
+ m1_n33990_17300# m1_n33750_9350# VSUBS VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt_WA2NKZ
XXM13 VSUBS m1_n30380_9040# m4_n15170_4960# VSUBS m1_n30380_9040# m4_n15170_4960#
+ sky130_fd_pr__nfet_01v8_lvt_QW8YAA
XXM37 m1_n37110_25500# m1_n41520_15180# m1_n37110_25500# m1_n35870_27710# m1_n41520_15180#
+ m1_n35870_27710# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_MXC9RL
Xsky130_fd_pr__nfet_01v8_lvt_W9NHZX_0 m1_n37700_18110# VSUBS m1_n37960_16980# m1_n37390_17440#
+ sky130_fd_pr__nfet_01v8_lvt_W9NHZX
XXM26 m1_n41520_15180# m1_n41290_16950# m1_n41520_15180# m1_n41290_16950# w_n40780_17110#
+ w_n40780_17110# m1_n41520_15180# w_n40780_17110# sky130_fd_pr__pfet_01v8_M5XJZ4
Xsky130_fd_pr__nfet_01v8_lvt_W9NHZX_1 m1_n37960_16980# VSUBS m1_n37960_16980# m1_n37390_15270#
+ sky130_fd_pr__nfet_01v8_lvt_W9NHZX
XXM27 m1_n37960_16980# m1_n41520_15180# m1_n39200_16970# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_M7ZRRL
Xbias_generator_0 m1_n34620_8840# w_n40780_17110# VSUBS bias_generator
XXM16 m4_n15170_4960# m1_n34970_4340# m1_n34970_4340# m1_n40040_26330# m4_n15170_4960#
+ m1_n34970_4340# m1_n34970_4340# w_n40780_17110# m4_n15170_4960# m1_n40040_26330#
+ m4_n15170_4960# m4_n15170_4960# m1_n40040_26330# m1_n34970_4340# m1_n34970_4340#
+ m1_n40040_26330# m1_n34970_4340# m4_n15170_4960# m1_n34970_4340# m4_n15170_4960#
+ m1_n40040_26330# m1_n34970_4340# m1_n34970_4340# m1_n34970_4340# m1_n34970_4340#
+ m1_n40040_26330# m1_n34970_4340# m1_n34970_4340# m4_n15170_4960# m1_n34970_4340#
+ m1_n34970_4340# m1_n34970_4340# m4_n15170_4960# m1_n40040_26330# m1_n34970_4340#
+ m1_n34970_4340# m1_n34970_4340# m1_n34970_4340# m4_n15170_4960# m1_n40040_26330#
+ m4_n15170_4960# m1_n34970_4340# m1_n34970_4340# m4_n15170_4960# m1_n34970_4340#
+ m1_n34970_4340# m1_n34970_4340# m1_n40040_26330# m4_n15170_4960# m1_n40040_26330#
+ m4_n15170_4960# m1_n40040_26330# m4_n15170_4960# m1_n40040_26330# m1_n34970_4340#
+ m4_n15170_4960# m1_n40040_26330# m1_n40040_26330# m1_n40040_26330# m1_n34970_4340#
+ m4_n15170_4960# m1_n34970_4340# m1_n34970_4340# m1_n40040_26330# m1_n34970_4340#
+ m1_n34970_4340# sky130_fd_pr__pfet_01v8_lvt_545GKL
XXM17 m1_n37960_25540# m4_n35400_n620# VSUBS w_n40780_17110# sky130_fd_pr__pfet_01v8_M7ZEKL
Xsky130_fd_pr__nfet_01v8_lvt_C84B7J_0 m1_n36990_22880# VSUBS m1_n29270_20310# VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_C84B7J
XXM28 m1_n41520_15180# m1_n41520_15180# m1_n41290_16950# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_M7ZRRL
XXM18 m1_n37960_25540# m4_n15170_4960# VSUBS w_n40780_17110# sky130_fd_pr__pfet_01v8_M7ZEKL
Xsky130_fd_pr__nfet_01v8_lvt_SHAVFW_0 m1_n36990_22880# m1_n36990_22880# m4_n22010_n680#
+ m4_n22010_n680# m1_n36990_22880# m4_n22010_n680# VSUBS VSUBS m4_n22010_n680# m1_n36990_22880#
+ m4_n22010_n680# VSUBS m1_n36990_22880# m1_n36990_22880# m1_n36990_22880# m1_n36990_22880#
+ m1_n36990_22880# VSUBS VSUBS m1_n36990_22880# m4_n22010_n680# m1_n36990_22880# m1_n36990_22880#
+ m1_n36990_22880# VSUBS VSUBS m1_n36990_22880# m4_n22010_n680# m1_n36990_22880# m1_n36990_22880#
+ VSUBS VSUBS VSUBS VSUBS m1_n36990_22880# m1_n36990_22880# m1_n36990_22880# m4_n22010_n680#
+ VSUBS m1_n36990_22880# VSUBS VSUBS m1_n36990_22880# m1_n36990_22880# m1_n36990_22880#
+ m1_n36990_22880# m1_n36990_22880# VSUBS m4_n22010_n680# m4_n22010_n680# VSUBS VSUBS
+ m4_n22010_n680# m1_n36990_22880# VSUBS m1_n36990_22880# m1_n36990_22880# m4_n22010_n680#
+ VSUBS m4_n22010_n680# m4_n22010_n680# m1_n36990_22880# m1_n36990_22880# m4_n22010_n680#
+ m4_n22010_n680# m4_n22010_n680# m4_n22010_n680# m1_n36990_22880# m1_n36990_22880#
+ m1_n36990_22880# m1_n36990_22880# sky130_fd_pr__nfet_01v8_lvt_SHAVFW
XXM2 m4_n22010_n680# m4_n22010_n680# m4_n22010_n680# m1_n35870_27710# m1_n35870_27710#
+ m4_n22010_n680# m1_n35870_27710# w_n40780_17110# m1_n35870_27710# m4_n22010_n680#
+ m4_n22010_n680# m1_n35870_27710# m1_n35870_27710# m1_n35870_27710# m1_n35870_27710#
+ w_n40780_17110# m4_n22010_n680# m1_n35870_27710# m1_n35870_27710# m1_n35870_27710#
+ w_n40780_17110# w_n40780_17110# m4_n22010_n680# w_n40780_17110# m4_n22010_n680#
+ m1_n35870_27710# m1_n35870_27710# w_n40780_17110# m1_n35870_27710# w_n40780_17110#
+ m4_n22010_n680# w_n40780_17110# m4_n22010_n680# m1_n35870_27710# m1_n35870_27710#
+ w_n40780_17110# w_n40780_17110# m1_n35870_27710# m1_n35870_27710# m1_n35870_27710#
+ m1_n35870_27710# w_n40780_17110# w_n40780_17110# m1_n35870_27710# m1_n35870_27710#
+ m4_n22010_n680# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_QQJVLQ
Xsky130_fd_pr__pfet_01v8_MD8735_0 m1_n35020_25500# w_n40780_17110# m1_n35020_25500#
+ m1_n41520_15180# m1_n41520_15180# m1_n41520_15180# m1_n35020_25500# m1_n41520_15180#
+ w_n40780_17110# m1_n41520_15180# m1_n35020_25500# w_n40780_17110# m1_n41520_15180#
+ w_n40780_17110# w_n40780_17110# sky130_fd_pr__pfet_01v8_MD8735
Xsky130_fd_pr__nfet_01v8_lvt_WA2NKZ_0 m1_n34620_8840# m1_n34620_8840# m1_n34620_8840#
+ m1_n41520_15180# m1_n34620_8840# m1_n33990_17300# m1_n41520_15180# m1_n41520_15180#
+ m1_n41520_15180# m1_n41520_15180# m1_n34620_8840# m1_n33990_17300# m1_n33990_17300#
+ m1_n33990_17300# m1_n34620_8840# m1_n33990_17300# m1_n41520_15180# m1_n34620_8840#
+ m1_n34620_8840# VSUBS m1_n33990_17300# m1_n34620_8840# m1_n41520_15180# m1_n41520_15180#
+ m1_n33990_17300# m1_n41520_15180# m1_n41520_15180# m1_n34620_8840# m1_n33990_17300#
+ m1_n33990_17300# m1_n33990_17300# sky130_fd_pr__nfet_01v8_lvt_WA2NKZ
XXM4 m1_n31060_24310# VSUBS m1_n31060_24310# VSUBS sky130_fd_pr__nfet_01v8_lvt_Q53FMB
XXM5 m1_n35870_27710# VSUBS m1_n40050_29050# m1_n36990_22880# sky130_fd_pr__nfet_01v8_lvt_Q53FMB
XXM6 w_n40780_17110# m1_n31050_29000# m1_n31050_29000# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_PD3USF
XXM7 m1_n31050_29000# m1_n37700_18110# m1_n37700_18110# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_SLP2FE
Xsky130_fd_pr__pfet_01v8_MV5GT4_0 m1_n39200_19680# m1_n41520_15180# m1_n39200_19680#
+ w_n40780_17110# m1_n39200_19680# m1_n39200_19680# m1_n41520_15180# m1_n41520_15180#
+ m1_n41520_15180# m1_n41520_15180# m1_n39200_19680# m1_n41520_15180# m1_n41520_15180#
+ m1_n39200_19680# w_n40780_17110# w_n40780_17110# m1_n41520_15180# m1_n39200_19680#
+ w_n40780_17110# m1_n41520_15180# w_n40780_17110# w_n40780_17110# m1_n39200_19680#
+ m1_n41520_15180# m1_n41520_15180# m1_n41520_15180# w_n40780_17110# w_n40780_17110#
+ w_n40780_17110# sky130_fd_pr__pfet_01v8_MV5GT4
XXM8 m1_n35870_27710# m1_n37700_18110# m1_n36990_22880# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_SLP2FE
Xsky130_fd_pr__nfet_01v8_lvt_QW8YAA_0 VSUBS m1_n30380_9040# m4_n15170_4960# VSUBS
+ m1_n30380_9040# m4_n15170_4960# sky130_fd_pr__nfet_01v8_lvt_QW8YAA
Xsky130_fd_pr__nfet_01v8_lvt_QW8YAA_1 VSUBS m1_n30380_9040# m4_n35400_n620# VSUBS
+ m1_n30380_9040# m4_n35400_n620# sky130_fd_pr__nfet_01v8_lvt_QW8YAA
Xsky130_fd_pr__nfet_01v8_lvt_QW8YAA_2 VSUBS m1_n30380_9040# m1_n30380_9040# VSUBS
+ m1_n30380_9040# m1_n30380_9040# sky130_fd_pr__nfet_01v8_lvt_QW8YAA
XXC1 m1_n36990_22880# m4_n22010_n680# sky130_fd_pr__cap_mim_m3_1_A4BC7Z
XXC2 m1_n35870_27710# m4_n22010_n680# sky130_fd_pr__cap_mim_m3_1_A4BC7Z
Xsky130_fd_pr__nfet_01v8_lvt_Q53FMB_0 m1_n40050_29050# VSUBS m1_n40050_29050# m1_n31060_24310#
+ sky130_fd_pr__nfet_01v8_lvt_Q53FMB
Xsky130_fd_pr__pfet_01v8_lvt_545GKL_0 m4_n15170_4960# m1_n34970_4340# m1_n34970_4340#
+ m1_n40040_26330# m4_n15170_4960# m1_n34970_4340# m1_n34970_4340# w_n40780_17110#
+ m4_n15170_4960# m1_n40040_26330# m4_n15170_4960# m4_n15170_4960# m1_n40040_26330#
+ m1_n34970_4340# m1_n34970_4340# m1_n40040_26330# m1_n34970_4340# m4_n15170_4960#
+ m1_n34970_4340# m4_n15170_4960# m1_n40040_26330# m1_n34970_4340# m1_n34970_4340#
+ m1_n34970_4340# m1_n34970_4340# m1_n40040_26330# m1_n34970_4340# m1_n34970_4340#
+ m4_n15170_4960# m1_n34970_4340# m1_n34970_4340# m1_n34970_4340# m4_n15170_4960#
+ m1_n40040_26330# m1_n34970_4340# m1_n34970_4340# m1_n34970_4340# m1_n34970_4340#
+ m4_n15170_4960# m1_n40040_26330# m4_n15170_4960# m1_n34970_4340# m1_n34970_4340#
+ m4_n15170_4960# m1_n34970_4340# m1_n34970_4340# m1_n34970_4340# m1_n40040_26330#
+ m4_n15170_4960# m1_n40040_26330# m4_n15170_4960# m1_n40040_26330# m4_n15170_4960#
+ m1_n40040_26330# m1_n34970_4340# m4_n15170_4960# m1_n40040_26330# m1_n40040_26330#
+ m1_n40040_26330# m1_n34970_4340# m4_n15170_4960# m1_n34970_4340# m1_n34970_4340#
+ m1_n40040_26330# m1_n34970_4340# m1_n34970_4340# sky130_fd_pr__pfet_01v8_lvt_545GKL
Xsky130_fd_pr__pfet_01v8_lvt_MF6SRL_0 m1_n39200_19680# m1_n41520_15180# m1_n41520_15180#
+ m1_n39200_19680# m1_n39200_19680# m1_n39200_19680# m1_n37960_25540# m1_n37960_25540#
+ m1_n41520_15180# m1_n37960_25540# m1_n37960_25540# w_n40780_17110# m1_n41520_15180#
+ sky130_fd_pr__pfet_01v8_lvt_MF6SRL
Xsky130_fd_pr__pfet_01v8_lvt_545GKL_1 m4_n35400_n620# m1_n34970_n360# m1_n34970_n360#
+ m1_n40040_26330# m4_n35400_n620# m1_n34970_n360# m1_n34970_n360# w_n40780_17110#
+ m4_n35400_n620# m1_n40040_26330# m4_n35400_n620# m4_n35400_n620# m1_n40040_26330#
+ m1_n34970_n360# m1_n34970_n360# m1_n40040_26330# m1_n34970_n360# m4_n35400_n620#
+ m1_n34970_n360# m4_n35400_n620# m1_n40040_26330# m1_n34970_n360# m1_n34970_n360#
+ m1_n34970_n360# m1_n34970_n360# m1_n40040_26330# m1_n34970_n360# m1_n34970_n360#
+ m4_n35400_n620# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360# m4_n35400_n620#
+ m1_n40040_26330# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360#
+ m4_n35400_n620# m1_n40040_26330# m4_n35400_n620# m1_n34970_n360# m1_n34970_n360#
+ m4_n35400_n620# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360# m1_n40040_26330#
+ m4_n35400_n620# m1_n40040_26330# m4_n35400_n620# m1_n40040_26330# m4_n35400_n620#
+ m1_n40040_26330# m1_n34970_n360# m4_n35400_n620# m1_n40040_26330# m1_n40040_26330#
+ m1_n40040_26330# m1_n34970_n360# m4_n35400_n620# m1_n34970_n360# m1_n34970_n360#
+ m1_n40040_26330# m1_n34970_n360# m1_n34970_n360# sky130_fd_pr__pfet_01v8_lvt_545GKL
Xsky130_fd_pr__nfet_01v8_lvt_N28DAC_0 VSUBS m1_n33750_9350# VSUBS m1_n33750_9350#
+ sky130_fd_pr__nfet_01v8_lvt_N28DAC
XXC3 m4_n35400_n620# VSUBS sky130_fd_pr__cap_mim_m3_1_5HBWYY
Xsky130_fd_pr__pfet_01v8_M7ZEKL_0 m1_n22730_15510# VSUBS m1_n30380_9040# w_n40780_17110#
+ sky130_fd_pr__pfet_01v8_M7ZEKL
Xsky130_fd_pr__pfet_01v8_lvt_545GKL_2 m4_n35400_n620# m1_n34970_n360# m1_n34970_n360#
+ m1_n40040_26330# m4_n35400_n620# m1_n34970_n360# m1_n34970_n360# w_n40780_17110#
+ m4_n35400_n620# m1_n40040_26330# m4_n35400_n620# m4_n35400_n620# m1_n40040_26330#
+ m1_n34970_n360# m1_n34970_n360# m1_n40040_26330# m1_n34970_n360# m4_n35400_n620#
+ m1_n34970_n360# m4_n35400_n620# m1_n40040_26330# m1_n34970_n360# m1_n34970_n360#
+ m1_n34970_n360# m1_n34970_n360# m1_n40040_26330# m1_n34970_n360# m1_n34970_n360#
+ m4_n35400_n620# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360# m4_n35400_n620#
+ m1_n40040_26330# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360#
+ m4_n35400_n620# m1_n40040_26330# m4_n35400_n620# m1_n34970_n360# m1_n34970_n360#
+ m4_n35400_n620# m1_n34970_n360# m1_n34970_n360# m1_n34970_n360# m1_n40040_26330#
+ m4_n35400_n620# m1_n40040_26330# m4_n35400_n620# m1_n40040_26330# m4_n35400_n620#
+ m1_n40040_26330# m1_n34970_n360# m4_n35400_n620# m1_n40040_26330# m1_n40040_26330#
+ m1_n40040_26330# m1_n34970_n360# m4_n35400_n620# m1_n34970_n360# m1_n34970_n360#
+ m1_n40040_26330# m1_n34970_n360# m1_n34970_n360# sky130_fd_pr__pfet_01v8_lvt_545GKL
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_0 m4_n35400_n620# VSUBS sky130_fd_pr__cap_mim_m3_1_5HBWYY
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_1 m4_n35400_n620# VSUBS sky130_fd_pr__cap_mim_m3_1_5HBWYY
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_2 m4_n35400_n620# VSUBS sky130_fd_pr__cap_mim_m3_1_5HBWYY
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_3 m4_n15170_4960# m4_n22010_n680# sky130_fd_pr__cap_mim_m3_1_5HBWYY
XXM40 m1_n41290_19650# m1_n41520_15180# m1_n41290_19650# w_n40780_17110# m1_n41290_19650#
+ m1_n41290_19650# m1_n41520_15180# m1_n41520_15180# m1_n41520_15180# m1_n41520_15180#
+ m1_n41290_19650# m1_n41520_15180# m1_n41520_15180# m1_n41290_19650# w_n40780_17110#
+ w_n40780_17110# m1_n41520_15180# m1_n41290_19650# w_n40780_17110# m1_n41520_15180#
+ w_n40780_17110# w_n40780_17110# m1_n41290_19650# m1_n41520_15180# m1_n41520_15180#
+ m1_n41520_15180# w_n40780_17110# w_n40780_17110# w_n40780_17110# sky130_fd_pr__pfet_01v8_MV5GT4
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_4 m4_n15170_4960# m4_n22010_n680# sky130_fd_pr__cap_mim_m3_1_5HBWYY
Xsky130_fd_pr__pfet_01v8_JHT74A_0 m1_n36990_22880# w_n40780_17110# m4_n35400_n620#
+ m1_n36990_22880# m4_n35400_n620# m1_n33780_27710# sky130_fd_pr__pfet_01v8_JHT74A
XXM41 m1_n41290_19650# m1_n41520_15180# m1_n41520_15180# m1_n41290_19650# m1_n41290_19650#
+ m1_n41290_19650# m1_n40040_26330# m1_n40040_26330# m1_n41520_15180# m1_n40040_26330#
+ m1_n40040_26330# w_n40780_17110# m1_n41520_15180# sky130_fd_pr__pfet_01v8_lvt_MF6SRL
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_5 m4_n15170_4960# m4_n22010_n680# sky130_fd_pr__cap_mim_m3_1_5HBWYY
XXM31 m1_n37390_15270# VSUBS m1_n37390_15270# VSUBS sky130_fd_pr__nfet_01v8_lvt_FWQUH5
Xsky130_fd_pr__cap_mim_m3_1_5HBWYY_6 m4_n15170_4960# m4_n22010_n680# sky130_fd_pr__cap_mim_m3_1_5HBWYY
XXM10 VSUBS VSUBS m1_n29270_20310# m1_n29270_20310# sky130_fd_pr__nfet_01v8_lvt_C84B7J
XXM21 VSUBS m1_n34620_8840# m1_n33750_9350# m1_n34620_8840# sky130_fd_pr__nfet_01v8_lvt_N28DAC
Xsky130_fd_pr__pfet_01v8_lvt_MXC9RL_0 m1_n35020_25500# m1_n41520_15180# m1_n35020_25500#
+ m1_n33780_27710# m1_n41520_15180# m1_n33780_27710# w_n40780_17110# sky130_fd_pr__pfet_01v8_lvt_MXC9RL
XXM44 m1_n37960_25540# m1_n22730_15510# w_n40780_17110# VSUBS sky130_fd_pr__pfet_01v8_F4HV3A
XXM11 m1_n29270_20310# w_n40780_17110# m4_n15170_4960# m1_n29270_20310# m4_n15170_4960#
+ m1_n33780_27710# sky130_fd_pr__pfet_01v8_JHT74A
Xsky130_fd_pr__nfet_01v8_lvt_FWQUH5_0 m1_n37390_17440# VSUBS m1_n37390_15270# VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_FWQUH5
.ends

