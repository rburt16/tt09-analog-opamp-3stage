magic
tech sky130A
magscale 1 2
timestamp 1730410385
<< pwell >>
rect -996 -279 996 279
<< nmos >>
rect -800 -131 800 69
<< ndiff >>
rect -858 57 -800 69
rect -858 -119 -846 57
rect -812 -119 -800 57
rect -858 -131 -800 -119
rect 800 57 858 69
rect 800 -119 812 57
rect 846 -119 858 57
rect 800 -131 858 -119
<< ndiffc >>
rect -846 -119 -812 57
rect 812 -119 846 57
<< psubdiff >>
rect -960 209 960 243
rect -960 -209 -926 209
rect 926 -209 960 209
rect -960 -243 -864 -209
rect 864 -243 960 -209
<< psubdiffcont >>
rect -864 -243 864 -209
<< poly >>
rect -800 141 800 157
rect -800 107 -784 141
rect 784 107 800 141
rect -800 69 800 107
rect -800 -157 800 -131
<< polycont >>
rect -784 107 784 141
<< locali >>
rect -960 209 960 243
rect -960 -209 -926 209
rect -800 107 -784 141
rect 784 107 800 141
rect -846 57 -812 73
rect -846 -135 -812 -119
rect 812 57 846 73
rect 812 -135 846 -119
rect 926 -209 960 209
rect -960 -243 -864 -209
rect 864 -243 960 -209
<< viali >>
rect -392 107 392 141
rect -846 -119 -812 57
rect 812 -119 846 57
rect -463 -243 463 -209
<< metal1 >>
rect -404 141 404 147
rect -404 107 -392 141
rect 392 107 404 141
rect -404 101 404 107
rect -852 57 -806 69
rect -852 -119 -846 57
rect -812 -119 -806 57
rect -852 -131 -806 -119
rect 806 57 852 69
rect 806 -119 812 57
rect 846 -119 852 57
rect 806 -131 852 -119
rect -475 -209 475 -203
rect -475 -243 -463 -209
rect 463 -243 475 -209
rect -475 -249 475 -243
<< properties >>
string FIXED_BBOX -943 -226 943 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 8.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 50 viagr 0 viagl 0 viagt 0
<< end >>
