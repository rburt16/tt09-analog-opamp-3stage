magic
tech sky130A
magscale 1 2
timestamp 1721946293
<< pwell >>
rect -1796 -221 1796 221
<< nmos >>
rect -1600 -73 1600 11
<< ndiff >>
rect -1658 -1 -1600 11
rect -1658 -61 -1646 -1
rect -1612 -61 -1600 -1
rect -1658 -73 -1600 -61
rect 1600 -1 1658 11
rect 1600 -61 1612 -1
rect 1646 -61 1658 -1
rect 1600 -73 1658 -61
<< ndiffc >>
rect -1646 -61 -1612 -1
rect 1612 -61 1646 -1
<< psubdiff >>
rect -1760 151 -1664 185
rect 1664 151 1760 185
rect -1760 89 -1726 151
rect 1726 89 1760 151
rect -1760 -151 -1726 -89
rect 1726 -151 1760 -89
rect -1760 -185 -1664 -151
rect 1664 -185 1760 -151
<< psubdiffcont >>
rect -1664 151 1664 185
rect -1760 -89 -1726 89
rect 1726 -89 1760 89
rect -1664 -185 1664 -151
<< poly >>
rect -1600 83 1600 99
rect -1600 49 -1584 83
rect 1584 49 1600 83
rect -1600 11 1600 49
rect -1600 -99 1600 -73
<< polycont >>
rect -1584 49 1584 83
<< locali >>
rect -1760 151 -1664 185
rect 1664 151 1760 185
rect -1760 89 -1726 151
rect 1726 89 1760 151
rect -1600 49 -1584 83
rect 1584 49 1600 83
rect -1646 -1 -1612 15
rect -1646 -77 -1612 -61
rect 1612 -1 1646 15
rect 1612 -77 1646 -61
rect -1760 -151 -1726 -89
rect 1726 -151 1760 -89
rect -1760 -185 -1664 -151
rect 1664 -185 1760 -151
<< viali >>
rect -792 49 792 83
rect -1646 -61 -1612 -1
rect 1612 -61 1646 -1
<< metal1 >>
rect -804 83 804 89
rect -804 49 -792 83
rect 792 49 804 83
rect -804 43 804 49
rect -1652 -1 -1606 11
rect -1652 -61 -1646 -1
rect -1612 -61 -1606 -1
rect -1652 -73 -1606 -61
rect 1606 -1 1652 11
rect 1606 -61 1612 -1
rect 1646 -61 1652 -1
rect 1606 -73 1652 -61
<< properties >>
string FIXED_BBOX -1743 -168 1743 168
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 16.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
