magic
tech sky130A
magscale 1 2
timestamp 1730482424
<< pwell >>
rect -596 -1010 596 1010
<< nmoslvt >>
rect -400 -800 400 800
<< ndiff >>
rect -458 552 -400 800
rect -458 -552 -446 552
rect -412 -552 -400 552
rect -458 -800 -400 -552
rect 400 552 458 800
rect 400 -552 412 552
rect 446 -552 458 552
rect 400 -800 458 -552
<< ndiffc >>
rect -446 -552 -412 552
rect 412 -552 446 552
<< psubdiff >>
rect -560 940 -325 974
rect 325 940 560 974
rect -560 615 -526 940
rect -560 -940 -526 -615
rect 526 615 560 940
rect 526 -940 560 -615
rect -560 -974 -325 -940
rect 325 -974 560 -940
<< psubdiffcont >>
rect -325 940 325 974
rect -560 -615 -526 615
rect 526 -615 560 615
rect -325 -974 325 -940
<< poly >>
rect -285 872 285 888
rect -285 855 -269 872
rect -400 838 -269 855
rect 269 855 285 872
rect 269 838 400 855
rect -400 800 400 838
rect -400 -838 400 -800
rect -400 -855 -269 -838
rect -285 -872 -269 -855
rect 269 -855 400 -838
rect 269 -872 285 -855
rect -285 -888 285 -872
<< polycont >>
rect -269 838 269 872
rect -269 -872 269 -838
<< locali >>
rect -560 940 -368 974
rect 368 940 560 974
rect -560 658 -526 940
rect 526 658 560 940
rect -446 552 -412 568
rect -446 -568 -412 -552
rect 412 552 446 568
rect 412 -568 446 -552
rect -560 -940 -526 -658
rect 526 -940 560 -658
rect -560 -974 -368 -940
rect 368 -974 560 -940
<< viali >>
rect -368 940 -325 974
rect -325 940 325 974
rect 325 940 368 974
rect -384 838 -269 872
rect -269 838 269 872
rect 269 838 384 872
rect -560 615 -526 658
rect -560 -615 -526 615
rect 526 615 560 658
rect -446 -552 -412 552
rect 412 -552 446 552
rect -560 -658 -526 -615
rect 526 -615 560 615
rect 526 -658 560 -615
rect -384 -872 -269 -838
rect -269 -872 269 -838
rect 269 -872 384 -838
rect -368 -974 -325 -940
rect -325 -974 325 -940
rect 325 -974 368 -940
<< metal1 >>
rect -380 974 380 980
rect -380 940 -368 974
rect 368 940 380 974
rect -380 934 380 940
rect -396 872 396 878
rect -396 838 -384 872
rect 384 838 396 872
rect -396 832 396 838
rect -566 658 -520 670
rect -566 -658 -560 658
rect -526 -658 -520 658
rect 520 658 566 670
rect -452 552 -406 564
rect -452 -552 -446 552
rect -412 -552 -406 552
rect -452 -564 -406 -552
rect 406 552 452 564
rect 406 -552 412 552
rect 446 -552 452 552
rect 406 -564 452 -552
rect -566 -670 -520 -658
rect 520 -658 526 658
rect 560 -658 566 658
rect 520 -670 566 -658
rect -396 -838 396 -832
rect -396 -872 -384 -838
rect 384 -872 396 -838
rect -396 -878 396 -872
rect -380 -940 380 -934
rect -380 -974 -368 -940
rect 368 -974 380 -940
rect -380 -980 380 -974
<< properties >>
string FIXED_BBOX -543 -957 543 957
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8.0 l 4.0 m 1 nf 1 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
