magic
tech sky130A
magscale 1 2
timestamp 1729896963
<< error_p >>
rect -1055 681 -993 687
rect -927 681 -865 687
rect -799 681 -737 687
rect -671 681 -609 687
rect -543 681 -481 687
rect -415 681 -353 687
rect -287 681 -225 687
rect -159 681 -97 687
rect -31 681 31 687
rect 97 681 159 687
rect 225 681 287 687
rect 353 681 415 687
rect 481 681 543 687
rect 609 681 671 687
rect 737 681 799 687
rect 865 681 927 687
rect 993 681 1055 687
rect -1055 647 -1043 681
rect -927 647 -915 681
rect -799 647 -787 681
rect -671 647 -659 681
rect -543 647 -531 681
rect -415 647 -403 681
rect -287 647 -275 681
rect -159 647 -147 681
rect -31 647 -19 681
rect 97 647 109 681
rect 225 647 237 681
rect 353 647 365 681
rect 481 647 493 681
rect 609 647 621 681
rect 737 647 749 681
rect 865 647 877 681
rect 993 647 1005 681
rect -1055 641 -993 647
rect -927 641 -865 647
rect -799 641 -737 647
rect -671 641 -609 647
rect -543 641 -481 647
rect -415 641 -353 647
rect -287 641 -225 647
rect -159 641 -97 647
rect -31 641 31 647
rect 97 641 159 647
rect 225 641 287 647
rect 353 641 415 647
rect 481 641 543 647
rect 609 641 671 647
rect 737 641 799 647
rect 865 641 927 647
rect 993 641 1055 647
rect -1055 71 -993 77
rect -927 71 -865 77
rect -799 71 -737 77
rect -671 71 -609 77
rect -543 71 -481 77
rect -415 71 -353 77
rect -287 71 -225 77
rect -159 71 -97 77
rect -31 71 31 77
rect 97 71 159 77
rect 225 71 287 77
rect 353 71 415 77
rect 481 71 543 77
rect 609 71 671 77
rect 737 71 799 77
rect 865 71 927 77
rect 993 71 1055 77
rect -1055 37 -1043 71
rect -927 37 -915 71
rect -799 37 -787 71
rect -671 37 -659 71
rect -543 37 -531 71
rect -415 37 -403 71
rect -287 37 -275 71
rect -159 37 -147 71
rect -31 37 -19 71
rect 97 37 109 71
rect 225 37 237 71
rect 353 37 365 71
rect 481 37 493 71
rect 609 37 621 71
rect 737 37 749 71
rect 865 37 877 71
rect 993 37 1005 71
rect -1055 31 -993 37
rect -927 31 -865 37
rect -799 31 -737 37
rect -671 31 -609 37
rect -543 31 -481 37
rect -415 31 -353 37
rect -287 31 -225 37
rect -159 31 -97 37
rect -31 31 31 37
rect 97 31 159 37
rect 225 31 287 37
rect 353 31 415 37
rect 481 31 543 37
rect 609 31 671 37
rect 737 31 799 37
rect 865 31 927 37
rect 993 31 1055 37
rect -1055 -37 -993 -31
rect -927 -37 -865 -31
rect -799 -37 -737 -31
rect -671 -37 -609 -31
rect -543 -37 -481 -31
rect -415 -37 -353 -31
rect -287 -37 -225 -31
rect -159 -37 -97 -31
rect -31 -37 31 -31
rect 97 -37 159 -31
rect 225 -37 287 -31
rect 353 -37 415 -31
rect 481 -37 543 -31
rect 609 -37 671 -31
rect 737 -37 799 -31
rect 865 -37 927 -31
rect 993 -37 1055 -31
rect -1055 -71 -1043 -37
rect -927 -71 -915 -37
rect -799 -71 -787 -37
rect -671 -71 -659 -37
rect -543 -71 -531 -37
rect -415 -71 -403 -37
rect -287 -71 -275 -37
rect -159 -71 -147 -37
rect -31 -71 -19 -37
rect 97 -71 109 -37
rect 225 -71 237 -37
rect 353 -71 365 -37
rect 481 -71 493 -37
rect 609 -71 621 -37
rect 737 -71 749 -37
rect 865 -71 877 -37
rect 993 -71 1005 -37
rect -1055 -77 -993 -71
rect -927 -77 -865 -71
rect -799 -77 -737 -71
rect -671 -77 -609 -71
rect -543 -77 -481 -71
rect -415 -77 -353 -71
rect -287 -77 -225 -71
rect -159 -77 -97 -71
rect -31 -77 31 -71
rect 97 -77 159 -71
rect 225 -77 287 -71
rect 353 -77 415 -71
rect 481 -77 543 -71
rect 609 -77 671 -71
rect 737 -77 799 -71
rect 865 -77 927 -71
rect 993 -77 1055 -71
rect -1055 -647 -993 -641
rect -927 -647 -865 -641
rect -799 -647 -737 -641
rect -671 -647 -609 -641
rect -543 -647 -481 -641
rect -415 -647 -353 -641
rect -287 -647 -225 -641
rect -159 -647 -97 -641
rect -31 -647 31 -641
rect 97 -647 159 -641
rect 225 -647 287 -641
rect 353 -647 415 -641
rect 481 -647 543 -641
rect 609 -647 671 -641
rect 737 -647 799 -641
rect 865 -647 927 -641
rect 993 -647 1055 -641
rect -1055 -681 -1043 -647
rect -927 -681 -915 -647
rect -799 -681 -787 -647
rect -671 -681 -659 -647
rect -543 -681 -531 -647
rect -415 -681 -403 -647
rect -287 -681 -275 -647
rect -159 -681 -147 -647
rect -31 -681 -19 -647
rect 97 -681 109 -647
rect 225 -681 237 -647
rect 353 -681 365 -647
rect 481 -681 493 -647
rect 609 -681 621 -647
rect 737 -681 749 -647
rect 865 -681 877 -647
rect 993 -681 1005 -647
rect -1055 -687 -993 -681
rect -927 -687 -865 -681
rect -799 -687 -737 -681
rect -671 -687 -609 -681
rect -543 -687 -481 -681
rect -415 -687 -353 -681
rect -287 -687 -225 -681
rect -159 -687 -97 -681
rect -31 -687 31 -681
rect 97 -687 159 -681
rect 225 -687 287 -681
rect 353 -687 415 -681
rect 481 -687 543 -681
rect 609 -687 671 -681
rect 737 -687 799 -681
rect 865 -687 927 -681
rect 993 -687 1055 -681
<< pwell >>
rect -1255 -819 1255 819
<< nmoslvt >>
rect -1059 109 -989 609
rect -931 109 -861 609
rect -803 109 -733 609
rect -675 109 -605 609
rect -547 109 -477 609
rect -419 109 -349 609
rect -291 109 -221 609
rect -163 109 -93 609
rect -35 109 35 609
rect 93 109 163 609
rect 221 109 291 609
rect 349 109 419 609
rect 477 109 547 609
rect 605 109 675 609
rect 733 109 803 609
rect 861 109 931 609
rect 989 109 1059 609
rect -1059 -609 -989 -109
rect -931 -609 -861 -109
rect -803 -609 -733 -109
rect -675 -609 -605 -109
rect -547 -609 -477 -109
rect -419 -609 -349 -109
rect -291 -609 -221 -109
rect -163 -609 -93 -109
rect -35 -609 35 -109
rect 93 -609 163 -109
rect 221 -609 291 -109
rect 349 -609 419 -109
rect 477 -609 547 -109
rect 605 -609 675 -109
rect 733 -609 803 -109
rect 861 -609 931 -109
rect 989 -609 1059 -109
<< ndiff >>
rect -1117 478 -1059 609
rect -1117 240 -1105 478
rect -1071 240 -1059 478
rect -1117 109 -1059 240
rect -989 478 -931 609
rect -989 240 -977 478
rect -943 240 -931 478
rect -989 109 -931 240
rect -861 478 -803 609
rect -861 240 -849 478
rect -815 240 -803 478
rect -861 109 -803 240
rect -733 478 -675 609
rect -733 240 -721 478
rect -687 240 -675 478
rect -733 109 -675 240
rect -605 478 -547 609
rect -605 240 -593 478
rect -559 240 -547 478
rect -605 109 -547 240
rect -477 478 -419 609
rect -477 240 -465 478
rect -431 240 -419 478
rect -477 109 -419 240
rect -349 478 -291 609
rect -349 240 -337 478
rect -303 240 -291 478
rect -349 109 -291 240
rect -221 478 -163 609
rect -221 240 -209 478
rect -175 240 -163 478
rect -221 109 -163 240
rect -93 478 -35 609
rect -93 240 -81 478
rect -47 240 -35 478
rect -93 109 -35 240
rect 35 478 93 609
rect 35 240 47 478
rect 81 240 93 478
rect 35 109 93 240
rect 163 478 221 609
rect 163 240 175 478
rect 209 240 221 478
rect 163 109 221 240
rect 291 478 349 609
rect 291 240 303 478
rect 337 240 349 478
rect 291 109 349 240
rect 419 478 477 609
rect 419 240 431 478
rect 465 240 477 478
rect 419 109 477 240
rect 547 478 605 609
rect 547 240 559 478
rect 593 240 605 478
rect 547 109 605 240
rect 675 478 733 609
rect 675 240 687 478
rect 721 240 733 478
rect 675 109 733 240
rect 803 478 861 609
rect 803 240 815 478
rect 849 240 861 478
rect 803 109 861 240
rect 931 478 989 609
rect 931 240 943 478
rect 977 240 989 478
rect 931 109 989 240
rect 1059 478 1117 609
rect 1059 240 1071 478
rect 1105 240 1117 478
rect 1059 109 1117 240
rect -1117 -240 -1059 -109
rect -1117 -478 -1105 -240
rect -1071 -478 -1059 -240
rect -1117 -609 -1059 -478
rect -989 -240 -931 -109
rect -989 -478 -977 -240
rect -943 -478 -931 -240
rect -989 -609 -931 -478
rect -861 -240 -803 -109
rect -861 -478 -849 -240
rect -815 -478 -803 -240
rect -861 -609 -803 -478
rect -733 -240 -675 -109
rect -733 -478 -721 -240
rect -687 -478 -675 -240
rect -733 -609 -675 -478
rect -605 -240 -547 -109
rect -605 -478 -593 -240
rect -559 -478 -547 -240
rect -605 -609 -547 -478
rect -477 -240 -419 -109
rect -477 -478 -465 -240
rect -431 -478 -419 -240
rect -477 -609 -419 -478
rect -349 -240 -291 -109
rect -349 -478 -337 -240
rect -303 -478 -291 -240
rect -349 -609 -291 -478
rect -221 -240 -163 -109
rect -221 -478 -209 -240
rect -175 -478 -163 -240
rect -221 -609 -163 -478
rect -93 -240 -35 -109
rect -93 -478 -81 -240
rect -47 -478 -35 -240
rect -93 -609 -35 -478
rect 35 -240 93 -109
rect 35 -478 47 -240
rect 81 -478 93 -240
rect 35 -609 93 -478
rect 163 -240 221 -109
rect 163 -478 175 -240
rect 209 -478 221 -240
rect 163 -609 221 -478
rect 291 -240 349 -109
rect 291 -478 303 -240
rect 337 -478 349 -240
rect 291 -609 349 -478
rect 419 -240 477 -109
rect 419 -478 431 -240
rect 465 -478 477 -240
rect 419 -609 477 -478
rect 547 -240 605 -109
rect 547 -478 559 -240
rect 593 -478 605 -240
rect 547 -609 605 -478
rect 675 -240 733 -109
rect 675 -478 687 -240
rect 721 -478 733 -240
rect 675 -609 733 -478
rect 803 -240 861 -109
rect 803 -478 815 -240
rect 849 -478 861 -240
rect 803 -609 861 -478
rect 931 -240 989 -109
rect 931 -478 943 -240
rect 977 -478 989 -240
rect 931 -609 989 -478
rect 1059 -240 1117 -109
rect 1059 -478 1071 -240
rect 1105 -478 1117 -240
rect 1059 -609 1117 -478
<< ndiffc >>
rect -1105 240 -1071 478
rect -977 240 -943 478
rect -849 240 -815 478
rect -721 240 -687 478
rect -593 240 -559 478
rect -465 240 -431 478
rect -337 240 -303 478
rect -209 240 -175 478
rect -81 240 -47 478
rect 47 240 81 478
rect 175 240 209 478
rect 303 240 337 478
rect 431 240 465 478
rect 559 240 593 478
rect 687 240 721 478
rect 815 240 849 478
rect 943 240 977 478
rect 1071 240 1105 478
rect -1105 -478 -1071 -240
rect -977 -478 -943 -240
rect -849 -478 -815 -240
rect -721 -478 -687 -240
rect -593 -478 -559 -240
rect -465 -478 -431 -240
rect -337 -478 -303 -240
rect -209 -478 -175 -240
rect -81 -478 -47 -240
rect 47 -478 81 -240
rect 175 -478 209 -240
rect 303 -478 337 -240
rect 431 -478 465 -240
rect 559 -478 593 -240
rect 687 -478 721 -240
rect 815 -478 849 -240
rect 943 -478 977 -240
rect 1071 -478 1105 -240
<< psubdiff >>
rect -1219 749 1219 783
rect -1219 344 -1185 749
rect -1219 -749 -1185 -344
rect 1185 -749 1219 749
rect -1219 -783 1219 -749
<< psubdiffcont >>
rect -1219 -344 -1185 344
<< poly >>
rect -1057 681 -991 697
rect -1057 664 -1041 681
rect -1059 647 -1041 664
rect -1007 664 -991 681
rect -929 681 -863 697
rect -929 664 -913 681
rect -1007 647 -989 664
rect -1059 609 -989 647
rect -931 647 -913 664
rect -879 664 -863 681
rect -801 681 -735 697
rect -801 664 -785 681
rect -879 647 -861 664
rect -931 609 -861 647
rect -803 647 -785 664
rect -751 664 -735 681
rect -673 681 -607 697
rect -673 664 -657 681
rect -751 647 -733 664
rect -803 609 -733 647
rect -675 647 -657 664
rect -623 664 -607 681
rect -545 681 -479 697
rect -545 664 -529 681
rect -623 647 -605 664
rect -675 609 -605 647
rect -547 647 -529 664
rect -495 664 -479 681
rect -417 681 -351 697
rect -417 664 -401 681
rect -495 647 -477 664
rect -547 609 -477 647
rect -419 647 -401 664
rect -367 664 -351 681
rect -289 681 -223 697
rect -289 664 -273 681
rect -367 647 -349 664
rect -419 609 -349 647
rect -291 647 -273 664
rect -239 664 -223 681
rect -161 681 -95 697
rect -161 664 -145 681
rect -239 647 -221 664
rect -291 609 -221 647
rect -163 647 -145 664
rect -111 664 -95 681
rect -33 681 33 697
rect -33 664 -17 681
rect -111 647 -93 664
rect -163 609 -93 647
rect -35 647 -17 664
rect 17 664 33 681
rect 95 681 161 697
rect 95 664 111 681
rect 17 647 35 664
rect -35 609 35 647
rect 93 647 111 664
rect 145 664 161 681
rect 223 681 289 697
rect 223 664 239 681
rect 145 647 163 664
rect 93 609 163 647
rect 221 647 239 664
rect 273 664 289 681
rect 351 681 417 697
rect 351 664 367 681
rect 273 647 291 664
rect 221 609 291 647
rect 349 647 367 664
rect 401 664 417 681
rect 479 681 545 697
rect 479 664 495 681
rect 401 647 419 664
rect 349 609 419 647
rect 477 647 495 664
rect 529 664 545 681
rect 607 681 673 697
rect 607 664 623 681
rect 529 647 547 664
rect 477 609 547 647
rect 605 647 623 664
rect 657 664 673 681
rect 735 681 801 697
rect 735 664 751 681
rect 657 647 675 664
rect 605 609 675 647
rect 733 647 751 664
rect 785 664 801 681
rect 863 681 929 697
rect 863 664 879 681
rect 785 647 803 664
rect 733 609 803 647
rect 861 647 879 664
rect 913 664 929 681
rect 991 681 1057 697
rect 991 664 1007 681
rect 913 647 931 664
rect 861 609 931 647
rect 989 647 1007 664
rect 1041 664 1057 681
rect 1041 647 1059 664
rect 989 609 1059 647
rect -1059 71 -989 109
rect -1059 54 -1041 71
rect -1057 37 -1041 54
rect -1007 54 -989 71
rect -931 71 -861 109
rect -931 54 -913 71
rect -1007 37 -991 54
rect -1057 21 -991 37
rect -929 37 -913 54
rect -879 54 -861 71
rect -803 71 -733 109
rect -803 54 -785 71
rect -879 37 -863 54
rect -929 21 -863 37
rect -801 37 -785 54
rect -751 54 -733 71
rect -675 71 -605 109
rect -675 54 -657 71
rect -751 37 -735 54
rect -801 21 -735 37
rect -673 37 -657 54
rect -623 54 -605 71
rect -547 71 -477 109
rect -547 54 -529 71
rect -623 37 -607 54
rect -673 21 -607 37
rect -545 37 -529 54
rect -495 54 -477 71
rect -419 71 -349 109
rect -419 54 -401 71
rect -495 37 -479 54
rect -545 21 -479 37
rect -417 37 -401 54
rect -367 54 -349 71
rect -291 71 -221 109
rect -291 54 -273 71
rect -367 37 -351 54
rect -417 21 -351 37
rect -289 37 -273 54
rect -239 54 -221 71
rect -163 71 -93 109
rect -163 54 -145 71
rect -239 37 -223 54
rect -289 21 -223 37
rect -161 37 -145 54
rect -111 54 -93 71
rect -35 71 35 109
rect -35 54 -17 71
rect -111 37 -95 54
rect -161 21 -95 37
rect -33 37 -17 54
rect 17 54 35 71
rect 93 71 163 109
rect 93 54 111 71
rect 17 37 33 54
rect -33 21 33 37
rect 95 37 111 54
rect 145 54 163 71
rect 221 71 291 109
rect 221 54 239 71
rect 145 37 161 54
rect 95 21 161 37
rect 223 37 239 54
rect 273 54 291 71
rect 349 71 419 109
rect 349 54 367 71
rect 273 37 289 54
rect 223 21 289 37
rect 351 37 367 54
rect 401 54 419 71
rect 477 71 547 109
rect 477 54 495 71
rect 401 37 417 54
rect 351 21 417 37
rect 479 37 495 54
rect 529 54 547 71
rect 605 71 675 109
rect 605 54 623 71
rect 529 37 545 54
rect 479 21 545 37
rect 607 37 623 54
rect 657 54 675 71
rect 733 71 803 109
rect 733 54 751 71
rect 657 37 673 54
rect 607 21 673 37
rect 735 37 751 54
rect 785 54 803 71
rect 861 71 931 109
rect 861 54 879 71
rect 785 37 801 54
rect 735 21 801 37
rect 863 37 879 54
rect 913 54 931 71
rect 989 71 1059 109
rect 989 54 1007 71
rect 913 37 929 54
rect 863 21 929 37
rect 991 37 1007 54
rect 1041 54 1059 71
rect 1041 37 1057 54
rect 991 21 1057 37
rect -1057 -37 -991 -21
rect -1057 -54 -1041 -37
rect -1059 -71 -1041 -54
rect -1007 -54 -991 -37
rect -929 -37 -863 -21
rect -929 -54 -913 -37
rect -1007 -71 -989 -54
rect -1059 -109 -989 -71
rect -931 -71 -913 -54
rect -879 -54 -863 -37
rect -801 -37 -735 -21
rect -801 -54 -785 -37
rect -879 -71 -861 -54
rect -931 -109 -861 -71
rect -803 -71 -785 -54
rect -751 -54 -735 -37
rect -673 -37 -607 -21
rect -673 -54 -657 -37
rect -751 -71 -733 -54
rect -803 -109 -733 -71
rect -675 -71 -657 -54
rect -623 -54 -607 -37
rect -545 -37 -479 -21
rect -545 -54 -529 -37
rect -623 -71 -605 -54
rect -675 -109 -605 -71
rect -547 -71 -529 -54
rect -495 -54 -479 -37
rect -417 -37 -351 -21
rect -417 -54 -401 -37
rect -495 -71 -477 -54
rect -547 -109 -477 -71
rect -419 -71 -401 -54
rect -367 -54 -351 -37
rect -289 -37 -223 -21
rect -289 -54 -273 -37
rect -367 -71 -349 -54
rect -419 -109 -349 -71
rect -291 -71 -273 -54
rect -239 -54 -223 -37
rect -161 -37 -95 -21
rect -161 -54 -145 -37
rect -239 -71 -221 -54
rect -291 -109 -221 -71
rect -163 -71 -145 -54
rect -111 -54 -95 -37
rect -33 -37 33 -21
rect -33 -54 -17 -37
rect -111 -71 -93 -54
rect -163 -109 -93 -71
rect -35 -71 -17 -54
rect 17 -54 33 -37
rect 95 -37 161 -21
rect 95 -54 111 -37
rect 17 -71 35 -54
rect -35 -109 35 -71
rect 93 -71 111 -54
rect 145 -54 161 -37
rect 223 -37 289 -21
rect 223 -54 239 -37
rect 145 -71 163 -54
rect 93 -109 163 -71
rect 221 -71 239 -54
rect 273 -54 289 -37
rect 351 -37 417 -21
rect 351 -54 367 -37
rect 273 -71 291 -54
rect 221 -109 291 -71
rect 349 -71 367 -54
rect 401 -54 417 -37
rect 479 -37 545 -21
rect 479 -54 495 -37
rect 401 -71 419 -54
rect 349 -109 419 -71
rect 477 -71 495 -54
rect 529 -54 545 -37
rect 607 -37 673 -21
rect 607 -54 623 -37
rect 529 -71 547 -54
rect 477 -109 547 -71
rect 605 -71 623 -54
rect 657 -54 673 -37
rect 735 -37 801 -21
rect 735 -54 751 -37
rect 657 -71 675 -54
rect 605 -109 675 -71
rect 733 -71 751 -54
rect 785 -54 801 -37
rect 863 -37 929 -21
rect 863 -54 879 -37
rect 785 -71 803 -54
rect 733 -109 803 -71
rect 861 -71 879 -54
rect 913 -54 929 -37
rect 991 -37 1057 -21
rect 991 -54 1007 -37
rect 913 -71 931 -54
rect 861 -109 931 -71
rect 989 -71 1007 -54
rect 1041 -54 1057 -37
rect 1041 -71 1059 -54
rect 989 -109 1059 -71
rect -1059 -647 -989 -609
rect -1059 -664 -1041 -647
rect -1057 -681 -1041 -664
rect -1007 -664 -989 -647
rect -931 -647 -861 -609
rect -931 -664 -913 -647
rect -1007 -681 -991 -664
rect -1057 -697 -991 -681
rect -929 -681 -913 -664
rect -879 -664 -861 -647
rect -803 -647 -733 -609
rect -803 -664 -785 -647
rect -879 -681 -863 -664
rect -929 -697 -863 -681
rect -801 -681 -785 -664
rect -751 -664 -733 -647
rect -675 -647 -605 -609
rect -675 -664 -657 -647
rect -751 -681 -735 -664
rect -801 -697 -735 -681
rect -673 -681 -657 -664
rect -623 -664 -605 -647
rect -547 -647 -477 -609
rect -547 -664 -529 -647
rect -623 -681 -607 -664
rect -673 -697 -607 -681
rect -545 -681 -529 -664
rect -495 -664 -477 -647
rect -419 -647 -349 -609
rect -419 -664 -401 -647
rect -495 -681 -479 -664
rect -545 -697 -479 -681
rect -417 -681 -401 -664
rect -367 -664 -349 -647
rect -291 -647 -221 -609
rect -291 -664 -273 -647
rect -367 -681 -351 -664
rect -417 -697 -351 -681
rect -289 -681 -273 -664
rect -239 -664 -221 -647
rect -163 -647 -93 -609
rect -163 -664 -145 -647
rect -239 -681 -223 -664
rect -289 -697 -223 -681
rect -161 -681 -145 -664
rect -111 -664 -93 -647
rect -35 -647 35 -609
rect -35 -664 -17 -647
rect -111 -681 -95 -664
rect -161 -697 -95 -681
rect -33 -681 -17 -664
rect 17 -664 35 -647
rect 93 -647 163 -609
rect 93 -664 111 -647
rect 17 -681 33 -664
rect -33 -697 33 -681
rect 95 -681 111 -664
rect 145 -664 163 -647
rect 221 -647 291 -609
rect 221 -664 239 -647
rect 145 -681 161 -664
rect 95 -697 161 -681
rect 223 -681 239 -664
rect 273 -664 291 -647
rect 349 -647 419 -609
rect 349 -664 367 -647
rect 273 -681 289 -664
rect 223 -697 289 -681
rect 351 -681 367 -664
rect 401 -664 419 -647
rect 477 -647 547 -609
rect 477 -664 495 -647
rect 401 -681 417 -664
rect 351 -697 417 -681
rect 479 -681 495 -664
rect 529 -664 547 -647
rect 605 -647 675 -609
rect 605 -664 623 -647
rect 529 -681 545 -664
rect 479 -697 545 -681
rect 607 -681 623 -664
rect 657 -664 675 -647
rect 733 -647 803 -609
rect 733 -664 751 -647
rect 657 -681 673 -664
rect 607 -697 673 -681
rect 735 -681 751 -664
rect 785 -664 803 -647
rect 861 -647 931 -609
rect 861 -664 879 -647
rect 785 -681 801 -664
rect 735 -697 801 -681
rect 863 -681 879 -664
rect 913 -664 931 -647
rect 989 -647 1059 -609
rect 989 -664 1007 -647
rect 913 -681 929 -664
rect 863 -697 929 -681
rect 991 -681 1007 -664
rect 1041 -664 1059 -647
rect 1041 -681 1057 -664
rect 991 -697 1057 -681
<< polycont >>
rect -1041 647 -1007 681
rect -913 647 -879 681
rect -785 647 -751 681
rect -657 647 -623 681
rect -529 647 -495 681
rect -401 647 -367 681
rect -273 647 -239 681
rect -145 647 -111 681
rect -17 647 17 681
rect 111 647 145 681
rect 239 647 273 681
rect 367 647 401 681
rect 495 647 529 681
rect 623 647 657 681
rect 751 647 785 681
rect 879 647 913 681
rect 1007 647 1041 681
rect -1041 37 -1007 71
rect -913 37 -879 71
rect -785 37 -751 71
rect -657 37 -623 71
rect -529 37 -495 71
rect -401 37 -367 71
rect -273 37 -239 71
rect -145 37 -111 71
rect -17 37 17 71
rect 111 37 145 71
rect 239 37 273 71
rect 367 37 401 71
rect 495 37 529 71
rect 623 37 657 71
rect 751 37 785 71
rect 879 37 913 71
rect 1007 37 1041 71
rect -1041 -71 -1007 -37
rect -913 -71 -879 -37
rect -785 -71 -751 -37
rect -657 -71 -623 -37
rect -529 -71 -495 -37
rect -401 -71 -367 -37
rect -273 -71 -239 -37
rect -145 -71 -111 -37
rect -17 -71 17 -37
rect 111 -71 145 -37
rect 239 -71 273 -37
rect 367 -71 401 -37
rect 495 -71 529 -37
rect 623 -71 657 -37
rect 751 -71 785 -37
rect 879 -71 913 -37
rect 1007 -71 1041 -37
rect -1041 -681 -1007 -647
rect -913 -681 -879 -647
rect -785 -681 -751 -647
rect -657 -681 -623 -647
rect -529 -681 -495 -647
rect -401 -681 -367 -647
rect -273 -681 -239 -647
rect -145 -681 -111 -647
rect -17 -681 17 -647
rect 111 -681 145 -647
rect 239 -681 273 -647
rect 367 -681 401 -647
rect 495 -681 529 -647
rect 623 -681 657 -647
rect 751 -681 785 -647
rect 879 -681 913 -647
rect 1007 -681 1041 -647
<< locali >>
rect -1219 749 1219 783
rect -1219 375 -1185 749
rect -1057 647 -1043 681
rect -1005 647 -991 681
rect -929 647 -915 681
rect -877 647 -863 681
rect -801 647 -787 681
rect -749 647 -735 681
rect -673 647 -659 681
rect -621 647 -607 681
rect -545 647 -531 681
rect -493 647 -479 681
rect -417 647 -403 681
rect -365 647 -351 681
rect -289 647 -275 681
rect -237 647 -223 681
rect -161 647 -147 681
rect -109 647 -95 681
rect -33 647 -19 681
rect 19 647 33 681
rect 95 647 109 681
rect 147 647 161 681
rect 223 647 237 681
rect 275 647 289 681
rect 351 647 365 681
rect 403 647 417 681
rect 479 647 493 681
rect 531 647 545 681
rect 607 647 621 681
rect 659 647 673 681
rect 735 647 749 681
rect 787 647 801 681
rect 863 647 877 681
rect 915 647 929 681
rect 991 647 1005 681
rect 1043 647 1057 681
rect -1105 478 -1071 494
rect -1105 224 -1071 240
rect -977 478 -943 494
rect -977 224 -943 240
rect -849 478 -815 494
rect -849 224 -815 240
rect -721 478 -687 494
rect -721 224 -687 240
rect -593 478 -559 494
rect -593 224 -559 240
rect -465 478 -431 494
rect -465 224 -431 240
rect -337 478 -303 494
rect -337 224 -303 240
rect -209 478 -175 494
rect -209 224 -175 240
rect -81 478 -47 494
rect -81 224 -47 240
rect 47 478 81 494
rect 47 224 81 240
rect 175 478 209 494
rect 175 224 209 240
rect 303 478 337 494
rect 303 224 337 240
rect 431 478 465 494
rect 431 224 465 240
rect 559 478 593 494
rect 559 224 593 240
rect 687 478 721 494
rect 687 224 721 240
rect 815 478 849 494
rect 815 224 849 240
rect 943 478 977 494
rect 943 224 977 240
rect 1071 478 1105 494
rect 1071 224 1105 240
rect -1057 37 -1043 71
rect -1005 37 -991 71
rect -929 37 -915 71
rect -877 37 -863 71
rect -801 37 -787 71
rect -749 37 -735 71
rect -673 37 -659 71
rect -621 37 -607 71
rect -545 37 -531 71
rect -493 37 -479 71
rect -417 37 -403 71
rect -365 37 -351 71
rect -289 37 -275 71
rect -237 37 -223 71
rect -161 37 -147 71
rect -109 37 -95 71
rect -33 37 -19 71
rect 19 37 33 71
rect 95 37 109 71
rect 147 37 161 71
rect 223 37 237 71
rect 275 37 289 71
rect 351 37 365 71
rect 403 37 417 71
rect 479 37 493 71
rect 531 37 545 71
rect 607 37 621 71
rect 659 37 673 71
rect 735 37 749 71
rect 787 37 801 71
rect 863 37 877 71
rect 915 37 929 71
rect 991 37 1005 71
rect 1043 37 1057 71
rect -1057 -71 -1043 -37
rect -1005 -71 -991 -37
rect -929 -71 -915 -37
rect -877 -71 -863 -37
rect -801 -71 -787 -37
rect -749 -71 -735 -37
rect -673 -71 -659 -37
rect -621 -71 -607 -37
rect -545 -71 -531 -37
rect -493 -71 -479 -37
rect -417 -71 -403 -37
rect -365 -71 -351 -37
rect -289 -71 -275 -37
rect -237 -71 -223 -37
rect -161 -71 -147 -37
rect -109 -71 -95 -37
rect -33 -71 -19 -37
rect 19 -71 33 -37
rect 95 -71 109 -37
rect 147 -71 161 -37
rect 223 -71 237 -37
rect 275 -71 289 -37
rect 351 -71 365 -37
rect 403 -71 417 -37
rect 479 -71 493 -37
rect 531 -71 545 -37
rect 607 -71 621 -37
rect 659 -71 673 -37
rect 735 -71 749 -37
rect 787 -71 801 -37
rect 863 -71 877 -37
rect 915 -71 929 -37
rect 991 -71 1005 -37
rect 1043 -71 1057 -37
rect -1219 -749 -1185 -375
rect -1105 -240 -1071 -224
rect -1105 -494 -1071 -478
rect -977 -240 -943 -224
rect -977 -494 -943 -478
rect -849 -240 -815 -224
rect -849 -494 -815 -478
rect -721 -240 -687 -224
rect -721 -494 -687 -478
rect -593 -240 -559 -224
rect -593 -494 -559 -478
rect -465 -240 -431 -224
rect -465 -494 -431 -478
rect -337 -240 -303 -224
rect -337 -494 -303 -478
rect -209 -240 -175 -224
rect -209 -494 -175 -478
rect -81 -240 -47 -224
rect -81 -494 -47 -478
rect 47 -240 81 -224
rect 47 -494 81 -478
rect 175 -240 209 -224
rect 175 -494 209 -478
rect 303 -240 337 -224
rect 303 -494 337 -478
rect 431 -240 465 -224
rect 431 -494 465 -478
rect 559 -240 593 -224
rect 559 -494 593 -478
rect 687 -240 721 -224
rect 687 -494 721 -478
rect 815 -240 849 -224
rect 815 -494 849 -478
rect 943 -240 977 -224
rect 943 -494 977 -478
rect 1071 -240 1105 -224
rect 1071 -494 1105 -478
rect -1057 -681 -1043 -647
rect -1005 -681 -991 -647
rect -929 -681 -915 -647
rect -877 -681 -863 -647
rect -801 -681 -787 -647
rect -749 -681 -735 -647
rect -673 -681 -659 -647
rect -621 -681 -607 -647
rect -545 -681 -531 -647
rect -493 -681 -479 -647
rect -417 -681 -403 -647
rect -365 -681 -351 -647
rect -289 -681 -275 -647
rect -237 -681 -223 -647
rect -161 -681 -147 -647
rect -109 -681 -95 -647
rect -33 -681 -19 -647
rect 19 -681 33 -647
rect 95 -681 109 -647
rect 147 -681 161 -647
rect 223 -681 237 -647
rect 275 -681 289 -647
rect 351 -681 365 -647
rect 403 -681 417 -647
rect 479 -681 493 -647
rect 531 -681 545 -647
rect 607 -681 621 -647
rect 659 -681 673 -647
rect 735 -681 749 -647
rect 787 -681 801 -647
rect 863 -681 877 -647
rect 915 -681 929 -647
rect 991 -681 1005 -647
rect 1043 -681 1057 -647
rect 1185 -749 1219 749
rect -1219 -783 1219 -749
<< viali >>
rect -1043 647 -1041 681
rect -1041 647 -1007 681
rect -1007 647 -1005 681
rect -915 647 -913 681
rect -913 647 -879 681
rect -879 647 -877 681
rect -787 647 -785 681
rect -785 647 -751 681
rect -751 647 -749 681
rect -659 647 -657 681
rect -657 647 -623 681
rect -623 647 -621 681
rect -531 647 -529 681
rect -529 647 -495 681
rect -495 647 -493 681
rect -403 647 -401 681
rect -401 647 -367 681
rect -367 647 -365 681
rect -275 647 -273 681
rect -273 647 -239 681
rect -239 647 -237 681
rect -147 647 -145 681
rect -145 647 -111 681
rect -111 647 -109 681
rect -19 647 -17 681
rect -17 647 17 681
rect 17 647 19 681
rect 109 647 111 681
rect 111 647 145 681
rect 145 647 147 681
rect 237 647 239 681
rect 239 647 273 681
rect 273 647 275 681
rect 365 647 367 681
rect 367 647 401 681
rect 401 647 403 681
rect 493 647 495 681
rect 495 647 529 681
rect 529 647 531 681
rect 621 647 623 681
rect 623 647 657 681
rect 657 647 659 681
rect 749 647 751 681
rect 751 647 785 681
rect 785 647 787 681
rect 877 647 879 681
rect 879 647 913 681
rect 913 647 915 681
rect 1005 647 1007 681
rect 1007 647 1041 681
rect 1041 647 1043 681
rect -1219 344 -1185 375
rect -1219 -344 -1185 344
rect -1105 240 -1071 478
rect -977 240 -943 478
rect -849 240 -815 478
rect -721 240 -687 478
rect -593 240 -559 478
rect -465 240 -431 478
rect -337 240 -303 478
rect -209 240 -175 478
rect -81 240 -47 478
rect 47 240 81 478
rect 175 240 209 478
rect 303 240 337 478
rect 431 240 465 478
rect 559 240 593 478
rect 687 240 721 478
rect 815 240 849 478
rect 943 240 977 478
rect 1071 240 1105 478
rect -1043 37 -1041 71
rect -1041 37 -1007 71
rect -1007 37 -1005 71
rect -915 37 -913 71
rect -913 37 -879 71
rect -879 37 -877 71
rect -787 37 -785 71
rect -785 37 -751 71
rect -751 37 -749 71
rect -659 37 -657 71
rect -657 37 -623 71
rect -623 37 -621 71
rect -531 37 -529 71
rect -529 37 -495 71
rect -495 37 -493 71
rect -403 37 -401 71
rect -401 37 -367 71
rect -367 37 -365 71
rect -275 37 -273 71
rect -273 37 -239 71
rect -239 37 -237 71
rect -147 37 -145 71
rect -145 37 -111 71
rect -111 37 -109 71
rect -19 37 -17 71
rect -17 37 17 71
rect 17 37 19 71
rect 109 37 111 71
rect 111 37 145 71
rect 145 37 147 71
rect 237 37 239 71
rect 239 37 273 71
rect 273 37 275 71
rect 365 37 367 71
rect 367 37 401 71
rect 401 37 403 71
rect 493 37 495 71
rect 495 37 529 71
rect 529 37 531 71
rect 621 37 623 71
rect 623 37 657 71
rect 657 37 659 71
rect 749 37 751 71
rect 751 37 785 71
rect 785 37 787 71
rect 877 37 879 71
rect 879 37 913 71
rect 913 37 915 71
rect 1005 37 1007 71
rect 1007 37 1041 71
rect 1041 37 1043 71
rect -1043 -71 -1041 -37
rect -1041 -71 -1007 -37
rect -1007 -71 -1005 -37
rect -915 -71 -913 -37
rect -913 -71 -879 -37
rect -879 -71 -877 -37
rect -787 -71 -785 -37
rect -785 -71 -751 -37
rect -751 -71 -749 -37
rect -659 -71 -657 -37
rect -657 -71 -623 -37
rect -623 -71 -621 -37
rect -531 -71 -529 -37
rect -529 -71 -495 -37
rect -495 -71 -493 -37
rect -403 -71 -401 -37
rect -401 -71 -367 -37
rect -367 -71 -365 -37
rect -275 -71 -273 -37
rect -273 -71 -239 -37
rect -239 -71 -237 -37
rect -147 -71 -145 -37
rect -145 -71 -111 -37
rect -111 -71 -109 -37
rect -19 -71 -17 -37
rect -17 -71 17 -37
rect 17 -71 19 -37
rect 109 -71 111 -37
rect 111 -71 145 -37
rect 145 -71 147 -37
rect 237 -71 239 -37
rect 239 -71 273 -37
rect 273 -71 275 -37
rect 365 -71 367 -37
rect 367 -71 401 -37
rect 401 -71 403 -37
rect 493 -71 495 -37
rect 495 -71 529 -37
rect 529 -71 531 -37
rect 621 -71 623 -37
rect 623 -71 657 -37
rect 657 -71 659 -37
rect 749 -71 751 -37
rect 751 -71 785 -37
rect 785 -71 787 -37
rect 877 -71 879 -37
rect 879 -71 913 -37
rect 913 -71 915 -37
rect 1005 -71 1007 -37
rect 1007 -71 1041 -37
rect 1041 -71 1043 -37
rect -1219 -375 -1185 -344
rect -1105 -478 -1071 -240
rect -977 -478 -943 -240
rect -849 -478 -815 -240
rect -721 -478 -687 -240
rect -593 -478 -559 -240
rect -465 -478 -431 -240
rect -337 -478 -303 -240
rect -209 -478 -175 -240
rect -81 -478 -47 -240
rect 47 -478 81 -240
rect 175 -478 209 -240
rect 303 -478 337 -240
rect 431 -478 465 -240
rect 559 -478 593 -240
rect 687 -478 721 -240
rect 815 -478 849 -240
rect 943 -478 977 -240
rect 1071 -478 1105 -240
rect -1043 -681 -1041 -647
rect -1041 -681 -1007 -647
rect -1007 -681 -1005 -647
rect -915 -681 -913 -647
rect -913 -681 -879 -647
rect -879 -681 -877 -647
rect -787 -681 -785 -647
rect -785 -681 -751 -647
rect -751 -681 -749 -647
rect -659 -681 -657 -647
rect -657 -681 -623 -647
rect -623 -681 -621 -647
rect -531 -681 -529 -647
rect -529 -681 -495 -647
rect -495 -681 -493 -647
rect -403 -681 -401 -647
rect -401 -681 -367 -647
rect -367 -681 -365 -647
rect -275 -681 -273 -647
rect -273 -681 -239 -647
rect -239 -681 -237 -647
rect -147 -681 -145 -647
rect -145 -681 -111 -647
rect -111 -681 -109 -647
rect -19 -681 -17 -647
rect -17 -681 17 -647
rect 17 -681 19 -647
rect 109 -681 111 -647
rect 111 -681 145 -647
rect 145 -681 147 -647
rect 237 -681 239 -647
rect 239 -681 273 -647
rect 273 -681 275 -647
rect 365 -681 367 -647
rect 367 -681 401 -647
rect 401 -681 403 -647
rect 493 -681 495 -647
rect 495 -681 529 -647
rect 529 -681 531 -647
rect 621 -681 623 -647
rect 623 -681 657 -647
rect 657 -681 659 -647
rect 749 -681 751 -647
rect 751 -681 785 -647
rect 785 -681 787 -647
rect 877 -681 879 -647
rect 879 -681 913 -647
rect 913 -681 915 -647
rect 1005 -681 1007 -647
rect 1007 -681 1041 -647
rect 1041 -681 1043 -647
<< metal1 >>
rect -1055 681 -993 687
rect -1055 647 -1043 681
rect -1005 647 -993 681
rect -1055 641 -993 647
rect -927 681 -865 687
rect -927 647 -915 681
rect -877 647 -865 681
rect -927 641 -865 647
rect -799 681 -737 687
rect -799 647 -787 681
rect -749 647 -737 681
rect -799 641 -737 647
rect -671 681 -609 687
rect -671 647 -659 681
rect -621 647 -609 681
rect -671 641 -609 647
rect -543 681 -481 687
rect -543 647 -531 681
rect -493 647 -481 681
rect -543 641 -481 647
rect -415 681 -353 687
rect -415 647 -403 681
rect -365 647 -353 681
rect -415 641 -353 647
rect -287 681 -225 687
rect -287 647 -275 681
rect -237 647 -225 681
rect -287 641 -225 647
rect -159 681 -97 687
rect -159 647 -147 681
rect -109 647 -97 681
rect -159 641 -97 647
rect -31 681 31 687
rect -31 647 -19 681
rect 19 647 31 681
rect -31 641 31 647
rect 97 681 159 687
rect 97 647 109 681
rect 147 647 159 681
rect 97 641 159 647
rect 225 681 287 687
rect 225 647 237 681
rect 275 647 287 681
rect 225 641 287 647
rect 353 681 415 687
rect 353 647 365 681
rect 403 647 415 681
rect 353 641 415 647
rect 481 681 543 687
rect 481 647 493 681
rect 531 647 543 681
rect 481 641 543 647
rect 609 681 671 687
rect 609 647 621 681
rect 659 647 671 681
rect 609 641 671 647
rect 737 681 799 687
rect 737 647 749 681
rect 787 647 799 681
rect 737 641 799 647
rect 865 681 927 687
rect 865 647 877 681
rect 915 647 927 681
rect 865 641 927 647
rect 993 681 1055 687
rect 993 647 1005 681
rect 1043 647 1055 681
rect 993 641 1055 647
rect -1111 478 -1065 490
rect -1225 375 -1179 387
rect -1225 -375 -1219 375
rect -1185 -375 -1179 375
rect -1111 240 -1105 478
rect -1071 240 -1065 478
rect -1111 228 -1065 240
rect -983 478 -937 490
rect -983 240 -977 478
rect -943 240 -937 478
rect -983 228 -937 240
rect -855 478 -809 490
rect -855 240 -849 478
rect -815 240 -809 478
rect -855 228 -809 240
rect -727 478 -681 490
rect -727 240 -721 478
rect -687 240 -681 478
rect -727 228 -681 240
rect -599 478 -553 490
rect -599 240 -593 478
rect -559 240 -553 478
rect -599 228 -553 240
rect -471 478 -425 490
rect -471 240 -465 478
rect -431 240 -425 478
rect -471 228 -425 240
rect -343 478 -297 490
rect -343 240 -337 478
rect -303 240 -297 478
rect -343 228 -297 240
rect -215 478 -169 490
rect -215 240 -209 478
rect -175 240 -169 478
rect -215 228 -169 240
rect -87 478 -41 490
rect -87 240 -81 478
rect -47 240 -41 478
rect -87 228 -41 240
rect 41 478 87 490
rect 41 240 47 478
rect 81 240 87 478
rect 41 228 87 240
rect 169 478 215 490
rect 169 240 175 478
rect 209 240 215 478
rect 169 228 215 240
rect 297 478 343 490
rect 297 240 303 478
rect 337 240 343 478
rect 297 228 343 240
rect 425 478 471 490
rect 425 240 431 478
rect 465 240 471 478
rect 425 228 471 240
rect 553 478 599 490
rect 553 240 559 478
rect 593 240 599 478
rect 553 228 599 240
rect 681 478 727 490
rect 681 240 687 478
rect 721 240 727 478
rect 681 228 727 240
rect 809 478 855 490
rect 809 240 815 478
rect 849 240 855 478
rect 809 228 855 240
rect 937 478 983 490
rect 937 240 943 478
rect 977 240 983 478
rect 937 228 983 240
rect 1065 478 1111 490
rect 1065 240 1071 478
rect 1105 240 1111 478
rect 1065 228 1111 240
rect -1055 71 -993 77
rect -1055 37 -1043 71
rect -1005 37 -993 71
rect -1055 31 -993 37
rect -927 71 -865 77
rect -927 37 -915 71
rect -877 37 -865 71
rect -927 31 -865 37
rect -799 71 -737 77
rect -799 37 -787 71
rect -749 37 -737 71
rect -799 31 -737 37
rect -671 71 -609 77
rect -671 37 -659 71
rect -621 37 -609 71
rect -671 31 -609 37
rect -543 71 -481 77
rect -543 37 -531 71
rect -493 37 -481 71
rect -543 31 -481 37
rect -415 71 -353 77
rect -415 37 -403 71
rect -365 37 -353 71
rect -415 31 -353 37
rect -287 71 -225 77
rect -287 37 -275 71
rect -237 37 -225 71
rect -287 31 -225 37
rect -159 71 -97 77
rect -159 37 -147 71
rect -109 37 -97 71
rect -159 31 -97 37
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect 97 71 159 77
rect 97 37 109 71
rect 147 37 159 71
rect 97 31 159 37
rect 225 71 287 77
rect 225 37 237 71
rect 275 37 287 71
rect 225 31 287 37
rect 353 71 415 77
rect 353 37 365 71
rect 403 37 415 71
rect 353 31 415 37
rect 481 71 543 77
rect 481 37 493 71
rect 531 37 543 71
rect 481 31 543 37
rect 609 71 671 77
rect 609 37 621 71
rect 659 37 671 71
rect 609 31 671 37
rect 737 71 799 77
rect 737 37 749 71
rect 787 37 799 71
rect 737 31 799 37
rect 865 71 927 77
rect 865 37 877 71
rect 915 37 927 71
rect 865 31 927 37
rect 993 71 1055 77
rect 993 37 1005 71
rect 1043 37 1055 71
rect 993 31 1055 37
rect -1055 -37 -993 -31
rect -1055 -71 -1043 -37
rect -1005 -71 -993 -37
rect -1055 -77 -993 -71
rect -927 -37 -865 -31
rect -927 -71 -915 -37
rect -877 -71 -865 -37
rect -927 -77 -865 -71
rect -799 -37 -737 -31
rect -799 -71 -787 -37
rect -749 -71 -737 -37
rect -799 -77 -737 -71
rect -671 -37 -609 -31
rect -671 -71 -659 -37
rect -621 -71 -609 -37
rect -671 -77 -609 -71
rect -543 -37 -481 -31
rect -543 -71 -531 -37
rect -493 -71 -481 -37
rect -543 -77 -481 -71
rect -415 -37 -353 -31
rect -415 -71 -403 -37
rect -365 -71 -353 -37
rect -415 -77 -353 -71
rect -287 -37 -225 -31
rect -287 -71 -275 -37
rect -237 -71 -225 -37
rect -287 -77 -225 -71
rect -159 -37 -97 -31
rect -159 -71 -147 -37
rect -109 -71 -97 -37
rect -159 -77 -97 -71
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect 97 -37 159 -31
rect 97 -71 109 -37
rect 147 -71 159 -37
rect 97 -77 159 -71
rect 225 -37 287 -31
rect 225 -71 237 -37
rect 275 -71 287 -37
rect 225 -77 287 -71
rect 353 -37 415 -31
rect 353 -71 365 -37
rect 403 -71 415 -37
rect 353 -77 415 -71
rect 481 -37 543 -31
rect 481 -71 493 -37
rect 531 -71 543 -37
rect 481 -77 543 -71
rect 609 -37 671 -31
rect 609 -71 621 -37
rect 659 -71 671 -37
rect 609 -77 671 -71
rect 737 -37 799 -31
rect 737 -71 749 -37
rect 787 -71 799 -37
rect 737 -77 799 -71
rect 865 -37 927 -31
rect 865 -71 877 -37
rect 915 -71 927 -37
rect 865 -77 927 -71
rect 993 -37 1055 -31
rect 993 -71 1005 -37
rect 1043 -71 1055 -37
rect 993 -77 1055 -71
rect -1225 -387 -1179 -375
rect -1111 -240 -1065 -228
rect -1111 -478 -1105 -240
rect -1071 -478 -1065 -240
rect -1111 -490 -1065 -478
rect -983 -240 -937 -228
rect -983 -478 -977 -240
rect -943 -478 -937 -240
rect -983 -490 -937 -478
rect -855 -240 -809 -228
rect -855 -478 -849 -240
rect -815 -478 -809 -240
rect -855 -490 -809 -478
rect -727 -240 -681 -228
rect -727 -478 -721 -240
rect -687 -478 -681 -240
rect -727 -490 -681 -478
rect -599 -240 -553 -228
rect -599 -478 -593 -240
rect -559 -478 -553 -240
rect -599 -490 -553 -478
rect -471 -240 -425 -228
rect -471 -478 -465 -240
rect -431 -478 -425 -240
rect -471 -490 -425 -478
rect -343 -240 -297 -228
rect -343 -478 -337 -240
rect -303 -478 -297 -240
rect -343 -490 -297 -478
rect -215 -240 -169 -228
rect -215 -478 -209 -240
rect -175 -478 -169 -240
rect -215 -490 -169 -478
rect -87 -240 -41 -228
rect -87 -478 -81 -240
rect -47 -478 -41 -240
rect -87 -490 -41 -478
rect 41 -240 87 -228
rect 41 -478 47 -240
rect 81 -478 87 -240
rect 41 -490 87 -478
rect 169 -240 215 -228
rect 169 -478 175 -240
rect 209 -478 215 -240
rect 169 -490 215 -478
rect 297 -240 343 -228
rect 297 -478 303 -240
rect 337 -478 343 -240
rect 297 -490 343 -478
rect 425 -240 471 -228
rect 425 -478 431 -240
rect 465 -478 471 -240
rect 425 -490 471 -478
rect 553 -240 599 -228
rect 553 -478 559 -240
rect 593 -478 599 -240
rect 553 -490 599 -478
rect 681 -240 727 -228
rect 681 -478 687 -240
rect 721 -478 727 -240
rect 681 -490 727 -478
rect 809 -240 855 -228
rect 809 -478 815 -240
rect 849 -478 855 -240
rect 809 -490 855 -478
rect 937 -240 983 -228
rect 937 -478 943 -240
rect 977 -478 983 -240
rect 937 -490 983 -478
rect 1065 -240 1111 -228
rect 1065 -478 1071 -240
rect 1105 -478 1111 -240
rect 1065 -490 1111 -478
rect -1055 -647 -993 -641
rect -1055 -681 -1043 -647
rect -1005 -681 -993 -647
rect -1055 -687 -993 -681
rect -927 -647 -865 -641
rect -927 -681 -915 -647
rect -877 -681 -865 -647
rect -927 -687 -865 -681
rect -799 -647 -737 -641
rect -799 -681 -787 -647
rect -749 -681 -737 -647
rect -799 -687 -737 -681
rect -671 -647 -609 -641
rect -671 -681 -659 -647
rect -621 -681 -609 -647
rect -671 -687 -609 -681
rect -543 -647 -481 -641
rect -543 -681 -531 -647
rect -493 -681 -481 -647
rect -543 -687 -481 -681
rect -415 -647 -353 -641
rect -415 -681 -403 -647
rect -365 -681 -353 -647
rect -415 -687 -353 -681
rect -287 -647 -225 -641
rect -287 -681 -275 -647
rect -237 -681 -225 -647
rect -287 -687 -225 -681
rect -159 -647 -97 -641
rect -159 -681 -147 -647
rect -109 -681 -97 -647
rect -159 -687 -97 -681
rect -31 -647 31 -641
rect -31 -681 -19 -647
rect 19 -681 31 -647
rect -31 -687 31 -681
rect 97 -647 159 -641
rect 97 -681 109 -647
rect 147 -681 159 -647
rect 97 -687 159 -681
rect 225 -647 287 -641
rect 225 -681 237 -647
rect 275 -681 287 -647
rect 225 -687 287 -681
rect 353 -647 415 -641
rect 353 -681 365 -647
rect 403 -681 415 -647
rect 353 -687 415 -681
rect 481 -647 543 -641
rect 481 -681 493 -647
rect 531 -681 543 -647
rect 481 -687 543 -681
rect 609 -647 671 -641
rect 609 -681 621 -647
rect 659 -681 671 -647
rect 609 -687 671 -681
rect 737 -647 799 -641
rect 737 -681 749 -647
rect 787 -681 799 -647
rect 737 -687 799 -681
rect 865 -647 927 -641
rect 865 -681 877 -647
rect 915 -681 927 -647
rect 865 -687 927 -681
rect 993 -647 1055 -641
rect 993 -681 1005 -647
rect 1043 -681 1055 -647
rect 993 -687 1055 -681
<< properties >>
string FIXED_BBOX -1202 -766 1202 766
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.5 l 0.35 m 2 nf 17 diffcov 50 polycov 70 guard 1 glc 1 grc 0 gtc 0 gbc 0 tbcov 50 rlcov 50 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 50 viadrn 50 viagate 100 viagb 0 viagr 0 viagl 50 viagt 0
<< end >>
