magic
tech sky130A
magscale 1 2
timestamp 1730569394
<< pwell >>
rect -596 -1919 596 1919
<< nmoslvt >>
rect -400 109 400 1709
rect -400 -1709 400 -109
<< ndiff >>
rect -458 1461 -400 1709
rect -458 357 -446 1461
rect -412 357 -400 1461
rect -458 109 -400 357
rect 400 1461 458 1709
rect 400 357 412 1461
rect 446 357 458 1461
rect 400 109 458 357
rect -458 -357 -400 -109
rect -458 -1461 -446 -357
rect -412 -1461 -400 -357
rect -458 -1709 -400 -1461
rect 400 -357 458 -109
rect 400 -1461 412 -357
rect 446 -1461 458 -357
rect 400 -1709 458 -1461
<< ndiffc >>
rect -446 357 -412 1461
rect 412 357 446 1461
rect -446 -1461 -412 -357
rect 412 -1461 446 -357
<< psubdiff >>
rect -560 1849 -325 1883
rect 325 1849 560 1883
rect -560 1251 -526 1849
rect 526 1251 560 1849
rect -560 -1849 -526 -1251
rect 526 -1849 560 -1251
rect -560 -1883 -325 -1849
rect 325 -1883 560 -1849
<< psubdiffcont >>
rect -325 1849 325 1883
rect -560 -1251 -526 1251
rect 526 -1251 560 1251
rect -325 -1883 325 -1849
<< poly >>
rect -285 1781 285 1797
rect -285 1764 -269 1781
rect -400 1747 -269 1764
rect 269 1764 285 1781
rect 269 1747 400 1764
rect -400 1709 400 1747
rect -400 71 400 109
rect -400 54 -269 71
rect -285 37 -269 54
rect 269 54 400 71
rect 269 37 285 54
rect -285 21 285 37
rect -285 -37 285 -21
rect -285 -54 -269 -37
rect -400 -71 -269 -54
rect 269 -54 285 -37
rect 269 -71 400 -54
rect -400 -109 400 -71
rect -400 -1747 400 -1709
rect -400 -1764 -269 -1747
rect -285 -1781 -269 -1764
rect 269 -1764 400 -1747
rect 269 -1781 285 -1764
rect -285 -1797 285 -1781
<< polycont >>
rect -269 1747 269 1781
rect -269 37 269 71
rect -269 -71 269 -37
rect -269 -1781 269 -1747
<< locali >>
rect -560 1849 -368 1883
rect 368 1849 560 1883
rect -560 1294 -526 1849
rect -446 1461 -412 1477
rect -446 341 -412 357
rect 412 1461 446 1477
rect 412 341 446 357
rect 526 1294 560 1849
rect -560 -1849 -526 -1294
rect -446 -357 -412 -341
rect -446 -1477 -412 -1461
rect 412 -357 446 -341
rect 412 -1477 446 -1461
rect 526 -1849 560 -1294
rect -560 -1883 -368 -1849
rect 368 -1883 560 -1849
<< viali >>
rect -368 1849 -325 1883
rect -325 1849 325 1883
rect 325 1849 368 1883
rect -384 1747 -269 1781
rect -269 1747 269 1781
rect 269 1747 384 1781
rect -560 1251 -526 1294
rect -560 -1251 -526 1251
rect -446 357 -412 1461
rect 412 357 446 1461
rect 526 1251 560 1294
rect -384 37 -269 71
rect -269 37 269 71
rect 269 37 384 71
rect -384 -71 -269 -37
rect -269 -71 269 -37
rect 269 -71 384 -37
rect -560 -1294 -526 -1251
rect -446 -1461 -412 -357
rect 412 -1461 446 -357
rect 526 -1251 560 1251
rect 526 -1294 560 -1251
rect -384 -1781 -269 -1747
rect -269 -1781 269 -1747
rect 269 -1781 384 -1747
rect -368 -1883 -325 -1849
rect -325 -1883 325 -1849
rect 325 -1883 368 -1849
<< metal1 >>
rect -380 1883 380 1889
rect -380 1849 -368 1883
rect 368 1849 380 1883
rect -380 1843 380 1849
rect -396 1781 396 1787
rect -396 1747 -384 1781
rect 384 1747 396 1781
rect -396 1741 396 1747
rect -452 1461 -406 1473
rect -566 1294 -520 1306
rect -566 -1294 -560 1294
rect -526 -1294 -520 1294
rect -452 357 -446 1461
rect -412 357 -406 1461
rect -452 345 -406 357
rect 406 1461 452 1473
rect 406 357 412 1461
rect 446 357 452 1461
rect 406 345 452 357
rect 520 1294 566 1306
rect -396 71 396 77
rect -396 37 -384 71
rect 384 37 396 71
rect -396 31 396 37
rect -396 -37 396 -31
rect -396 -71 -384 -37
rect 384 -71 396 -37
rect -396 -77 396 -71
rect -566 -1306 -520 -1294
rect -452 -357 -406 -345
rect -452 -1461 -446 -357
rect -412 -1461 -406 -357
rect -452 -1473 -406 -1461
rect 406 -357 452 -345
rect 406 -1461 412 -357
rect 446 -1461 452 -357
rect 520 -1294 526 1294
rect 560 -1294 566 1294
rect 520 -1306 566 -1294
rect 406 -1473 452 -1461
rect -396 -1747 396 -1741
rect -396 -1781 -384 -1747
rect 384 -1781 396 -1747
rect -396 -1787 396 -1781
rect -380 -1849 380 -1843
rect -380 -1883 -368 -1849
rect 368 -1883 380 -1849
rect -380 -1889 380 -1883
<< properties >>
string FIXED_BBOX -543 -1866 543 1866
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 8.0 l 4.0 m 2 nf 1 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
