magic
tech sky130A
magscale 1 2
timestamp 1729617920
<< error_p >>
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect -31 2159 31 2165
rect -31 71 31 77
rect -31 37 -19 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect -31 -77 31 -71
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect -31 -2205 31 -2199
<< nwell >>
rect -231 -2337 231 2337
<< pmoslvt >>
rect -35 118 35 2118
rect -35 -2118 35 -118
<< pdiff >>
rect -93 2106 -35 2118
rect -93 130 -81 2106
rect -47 130 -35 2106
rect -93 118 -35 130
rect 35 2106 93 2118
rect 35 130 47 2106
rect 81 130 93 2106
rect 35 118 93 130
rect -93 -130 -35 -118
rect -93 -2106 -81 -130
rect -47 -2106 -35 -130
rect -93 -2118 -35 -2106
rect 35 -130 93 -118
rect 35 -2106 47 -130
rect 81 -2106 93 -130
rect 35 -2118 93 -2106
<< pdiffc >>
rect -81 130 -47 2106
rect 47 130 81 2106
rect -81 -2106 -47 -130
rect 47 -2106 81 -130
<< nsubdiff >>
rect -195 2267 -99 2301
rect 99 2267 195 2301
rect -195 2205 -161 2267
rect 161 2205 195 2267
rect -195 -2267 -161 -2205
rect 161 -2267 195 -2205
rect -195 -2301 -99 -2267
rect 99 -2301 195 -2267
<< nsubdiffcont >>
rect -99 2267 99 2301
rect -195 -2205 -161 2205
rect 161 -2205 195 2205
rect -99 -2301 99 -2267
<< poly >>
rect -35 2199 35 2215
rect -35 2165 -19 2199
rect 19 2165 35 2199
rect -35 2118 35 2165
rect -35 71 35 118
rect -35 37 -19 71
rect 19 37 35 71
rect -35 21 35 37
rect -35 -37 35 -21
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -35 -118 35 -71
rect -35 -2165 35 -2118
rect -35 -2199 -19 -2165
rect 19 -2199 35 -2165
rect -35 -2215 35 -2199
<< polycont >>
rect -19 2165 19 2199
rect -19 37 19 71
rect -19 -71 19 -37
rect -19 -2199 19 -2165
<< locali >>
rect -195 2267 -99 2301
rect 99 2267 195 2301
rect -195 2205 -161 2267
rect 161 2205 195 2267
rect -35 2165 -19 2199
rect 19 2165 35 2199
rect -81 2106 -47 2122
rect -81 114 -47 130
rect 47 2106 81 2122
rect 47 114 81 130
rect -35 37 -19 71
rect 19 37 35 71
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -81 -130 -47 -114
rect -81 -2122 -47 -2106
rect 47 -130 81 -114
rect 47 -2122 81 -2106
rect -35 -2199 -19 -2165
rect 19 -2199 35 -2165
rect -195 -2267 -161 -2205
rect 161 -2267 195 -2205
rect -195 -2301 -99 -2267
rect 99 -2301 195 -2267
<< viali >>
rect -19 2165 19 2199
rect -81 130 -47 2106
rect 47 130 81 2106
rect -19 37 19 71
rect -19 -71 19 -37
rect -81 -2106 -47 -130
rect 47 -2106 81 -130
rect -19 -2199 19 -2165
<< metal1 >>
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect 19 2165 31 2199
rect -31 2159 31 2165
rect -87 2106 -41 2118
rect -87 130 -81 2106
rect -47 130 -41 2106
rect -87 118 -41 130
rect 41 2106 87 2118
rect 41 130 47 2106
rect 81 130 87 2106
rect 41 118 87 130
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect -87 -130 -41 -118
rect -87 -2106 -81 -130
rect -47 -2106 -41 -130
rect -87 -2118 -41 -2106
rect 41 -130 87 -118
rect 41 -2106 47 -130
rect 81 -2106 87 -130
rect 41 -2118 87 -2106
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect 19 -2199 31 -2165
rect -31 -2205 31 -2199
<< properties >>
string FIXED_BBOX -178 -2284 178 2284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
