magic
tech sky130A
magscale 1 2
timestamp 1730569394
<< error_p >>
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect -31 2159 31 2165
rect -31 71 31 77
rect -31 37 -19 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect -31 -77 31 -71
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect -31 -2205 31 -2199
<< nwell >>
rect -231 -2337 231 2337
<< pmoslvt >>
rect -35 118 35 2118
rect -35 -2118 35 -118
<< pdiff >>
rect -93 1810 -35 2118
rect -93 426 -81 1810
rect -47 426 -35 1810
rect -93 118 -35 426
rect 35 1810 93 2118
rect 35 426 47 1810
rect 81 426 93 1810
rect 35 118 93 426
rect -93 -426 -35 -118
rect -93 -1810 -81 -426
rect -47 -1810 -35 -426
rect -93 -2118 -35 -1810
rect 35 -426 93 -118
rect 35 -1810 47 -426
rect 81 -1810 93 -426
rect 35 -2118 93 -1810
<< pdiffc >>
rect -81 426 -47 1810
rect 47 426 81 1810
rect -81 -1810 -47 -426
rect 47 -1810 81 -426
<< nsubdiff >>
rect -195 2267 -69 2301
rect 69 2267 195 2301
rect -195 1544 -161 2267
rect 161 1544 195 2267
rect -195 -2267 -161 -1544
rect 161 -2267 195 -1544
rect -195 -2301 -69 -2267
rect 69 -2301 195 -2267
<< nsubdiffcont >>
rect -69 2267 69 2301
rect -195 -1544 -161 1544
rect 161 -1544 195 1544
rect -69 -2301 69 -2267
<< poly >>
rect -33 2199 33 2215
rect -33 2182 -17 2199
rect -35 2165 -17 2182
rect 17 2182 33 2199
rect 17 2165 35 2182
rect -35 2118 35 2165
rect -35 71 35 118
rect -35 54 -17 71
rect -33 37 -17 54
rect 17 54 35 71
rect 17 37 33 54
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -54 -17 -37
rect -35 -71 -17 -54
rect 17 -54 33 -37
rect 17 -71 35 -54
rect -35 -118 35 -71
rect -35 -2165 35 -2118
rect -35 -2182 -17 -2165
rect -33 -2199 -17 -2182
rect 17 -2182 35 -2165
rect 17 -2199 33 -2182
rect -33 -2215 33 -2199
<< polycont >>
rect -17 2165 17 2199
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -2199 17 -2165
<< locali >>
rect -195 2267 -113 2301
rect 113 2267 195 2301
rect -195 1587 -161 2267
rect -33 2165 -19 2199
rect 19 2165 33 2199
rect -81 1810 -47 1826
rect -81 410 -47 426
rect 47 1810 81 1826
rect 47 410 81 426
rect 161 1587 195 2267
rect -33 37 -19 71
rect 19 37 33 71
rect -33 -71 -19 -37
rect 19 -71 33 -37
rect -195 -2267 -161 -1587
rect -81 -426 -47 -410
rect -81 -1826 -47 -1810
rect 47 -426 81 -410
rect 47 -1826 81 -1810
rect -33 -2199 -19 -2165
rect 19 -2199 33 -2165
rect 161 -2267 195 -1587
rect -195 -2301 -113 -2267
rect 113 -2301 195 -2267
<< viali >>
rect -113 2267 -69 2301
rect -69 2267 69 2301
rect 69 2267 113 2301
rect -19 2165 -17 2199
rect -17 2165 17 2199
rect 17 2165 19 2199
rect -195 1544 -161 1587
rect -195 -1544 -161 1544
rect -81 426 -47 1810
rect 47 426 81 1810
rect 161 1544 195 1587
rect -19 37 -17 71
rect -17 37 17 71
rect 17 37 19 71
rect -19 -71 -17 -37
rect -17 -71 17 -37
rect 17 -71 19 -37
rect -195 -1587 -161 -1544
rect -81 -1810 -47 -426
rect 47 -1810 81 -426
rect 161 -1544 195 1544
rect 161 -1587 195 -1544
rect -19 -2199 -17 -2165
rect -17 -2199 17 -2165
rect 17 -2199 19 -2165
rect -113 -2301 -69 -2267
rect -69 -2301 69 -2267
rect 69 -2301 113 -2267
<< metal1 >>
rect -125 2301 125 2307
rect -125 2267 -113 2301
rect 113 2267 125 2301
rect -125 2261 125 2267
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect 19 2165 31 2199
rect -31 2159 31 2165
rect -87 1810 -41 1822
rect -201 1587 -155 1599
rect -201 -1587 -195 1587
rect -161 -1587 -155 1587
rect -87 426 -81 1810
rect -47 426 -41 1810
rect -87 414 -41 426
rect 41 1810 87 1822
rect 41 426 47 1810
rect 81 426 87 1810
rect 41 414 87 426
rect 155 1587 201 1599
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect -201 -1599 -155 -1587
rect -87 -426 -41 -414
rect -87 -1810 -81 -426
rect -47 -1810 -41 -426
rect -87 -1822 -41 -1810
rect 41 -426 87 -414
rect 41 -1810 47 -426
rect 81 -1810 87 -426
rect 155 -1587 161 1587
rect 195 -1587 201 1587
rect 155 -1599 201 -1587
rect 41 -1822 87 -1810
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect 19 -2199 31 -2165
rect -31 -2205 31 -2199
rect -125 -2267 125 -2261
rect -125 -2301 -113 -2267
rect 113 -2301 125 -2267
rect -125 -2307 125 -2301
<< properties >>
string FIXED_BBOX -178 -2284 178 2284
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 2 nf 1 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
