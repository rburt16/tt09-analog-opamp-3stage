magic
tech sky130A
magscale 1 2
timestamp 1730482424
<< nwell >>
rect -554 -4573 554 4573
<< pmos >>
rect -358 2354 -158 4354
rect -100 2354 100 4354
rect 158 2354 358 4354
rect -358 118 -158 2118
rect -100 118 100 2118
rect 158 118 358 2118
rect -358 -2118 -158 -118
rect -100 -2118 100 -118
rect 158 -2118 358 -118
rect -358 -4354 -158 -2354
rect -100 -4354 100 -2354
rect 158 -4354 358 -2354
<< pdiff >>
rect -416 4046 -358 4354
rect -416 2662 -404 4046
rect -370 2662 -358 4046
rect -416 2354 -358 2662
rect -158 4046 -100 4354
rect -158 2662 -146 4046
rect -112 2662 -100 4046
rect -158 2354 -100 2662
rect 100 4046 158 4354
rect 100 2662 112 4046
rect 146 2662 158 4046
rect 100 2354 158 2662
rect 358 4046 416 4354
rect 358 2662 370 4046
rect 404 2662 416 4046
rect 358 2354 416 2662
rect -416 1810 -358 2118
rect -416 426 -404 1810
rect -370 426 -358 1810
rect -416 118 -358 426
rect -158 1810 -100 2118
rect -158 426 -146 1810
rect -112 426 -100 1810
rect -158 118 -100 426
rect 100 1810 158 2118
rect 100 426 112 1810
rect 146 426 158 1810
rect 100 118 158 426
rect 358 1810 416 2118
rect 358 426 370 1810
rect 404 426 416 1810
rect 358 118 416 426
rect -416 -426 -358 -118
rect -416 -1810 -404 -426
rect -370 -1810 -358 -426
rect -416 -2118 -358 -1810
rect -158 -426 -100 -118
rect -158 -1810 -146 -426
rect -112 -1810 -100 -426
rect -158 -2118 -100 -1810
rect 100 -426 158 -118
rect 100 -1810 112 -426
rect 146 -1810 158 -426
rect 100 -2118 158 -1810
rect 358 -426 416 -118
rect 358 -1810 370 -426
rect 404 -1810 416 -426
rect 358 -2118 416 -1810
rect -416 -2662 -358 -2354
rect -416 -4046 -404 -2662
rect -370 -4046 -358 -2662
rect -416 -4354 -358 -4046
rect -158 -2662 -100 -2354
rect -158 -4046 -146 -2662
rect -112 -4046 -100 -2662
rect -158 -4354 -100 -4046
rect 100 -2662 158 -2354
rect 100 -4046 112 -2662
rect 146 -4046 158 -2662
rect 100 -4354 158 -4046
rect 358 -2662 416 -2354
rect 358 -4046 370 -2662
rect 404 -4046 416 -2662
rect 358 -4354 416 -4046
<< pdiffc >>
rect -404 2662 -370 4046
rect -146 2662 -112 4046
rect 112 2662 146 4046
rect 370 2662 404 4046
rect -404 426 -370 1810
rect -146 426 -112 1810
rect 112 426 146 1810
rect 370 426 404 1810
rect -404 -1810 -370 -426
rect -146 -1810 -112 -426
rect 112 -1810 146 -426
rect 370 -1810 404 -426
rect -404 -4046 -370 -2662
rect -146 -4046 -112 -2662
rect 112 -4046 146 -2662
rect 370 -4046 404 -2662
<< nsubdiff >>
rect -518 4503 -295 4537
rect 295 4503 518 4537
rect -518 3109 -484 4503
rect 484 3109 518 4503
rect -518 -4503 -484 -3109
rect 484 -4503 518 -3109
rect -518 -4537 -295 -4503
rect 295 -4537 518 -4503
<< nsubdiffcont >>
rect -295 4503 295 4537
rect -518 -3109 -484 3109
rect 484 -3109 518 3109
rect -295 -4537 295 -4503
<< poly >>
rect -333 4435 -183 4451
rect -333 4418 -317 4435
rect -358 4401 -317 4418
rect -199 4418 -183 4435
rect -75 4435 75 4451
rect -75 4418 -59 4435
rect -199 4401 -158 4418
rect -358 4354 -158 4401
rect -100 4401 -59 4418
rect 59 4418 75 4435
rect 183 4435 333 4451
rect 183 4418 199 4435
rect 59 4401 100 4418
rect -100 4354 100 4401
rect 158 4401 199 4418
rect 317 4418 333 4435
rect 317 4401 358 4418
rect 158 4354 358 4401
rect -358 2307 -158 2354
rect -358 2290 -317 2307
rect -333 2273 -317 2290
rect -199 2290 -158 2307
rect -100 2307 100 2354
rect -100 2290 -59 2307
rect -199 2273 -183 2290
rect -333 2257 -183 2273
rect -75 2273 -59 2290
rect 59 2290 100 2307
rect 158 2307 358 2354
rect 158 2290 199 2307
rect 59 2273 75 2290
rect -75 2257 75 2273
rect 183 2273 199 2290
rect 317 2290 358 2307
rect 317 2273 333 2290
rect 183 2257 333 2273
rect -333 2199 -183 2215
rect -333 2182 -317 2199
rect -358 2165 -317 2182
rect -199 2182 -183 2199
rect -75 2199 75 2215
rect -75 2182 -59 2199
rect -199 2165 -158 2182
rect -358 2118 -158 2165
rect -100 2165 -59 2182
rect 59 2182 75 2199
rect 183 2199 333 2215
rect 183 2182 199 2199
rect 59 2165 100 2182
rect -100 2118 100 2165
rect 158 2165 199 2182
rect 317 2182 333 2199
rect 317 2165 358 2182
rect 158 2118 358 2165
rect -358 71 -158 118
rect -358 54 -317 71
rect -333 37 -317 54
rect -199 54 -158 71
rect -100 71 100 118
rect -100 54 -59 71
rect -199 37 -183 54
rect -333 21 -183 37
rect -75 37 -59 54
rect 59 54 100 71
rect 158 71 358 118
rect 158 54 199 71
rect 59 37 75 54
rect -75 21 75 37
rect 183 37 199 54
rect 317 54 358 71
rect 317 37 333 54
rect 183 21 333 37
rect -333 -37 -183 -21
rect -333 -54 -317 -37
rect -358 -71 -317 -54
rect -199 -54 -183 -37
rect -75 -37 75 -21
rect -75 -54 -59 -37
rect -199 -71 -158 -54
rect -358 -118 -158 -71
rect -100 -71 -59 -54
rect 59 -54 75 -37
rect 183 -37 333 -21
rect 183 -54 199 -37
rect 59 -71 100 -54
rect -100 -118 100 -71
rect 158 -71 199 -54
rect 317 -54 333 -37
rect 317 -71 358 -54
rect 158 -118 358 -71
rect -358 -2165 -158 -2118
rect -358 -2182 -317 -2165
rect -333 -2199 -317 -2182
rect -199 -2182 -158 -2165
rect -100 -2165 100 -2118
rect -100 -2182 -59 -2165
rect -199 -2199 -183 -2182
rect -333 -2215 -183 -2199
rect -75 -2199 -59 -2182
rect 59 -2182 100 -2165
rect 158 -2165 358 -2118
rect 158 -2182 199 -2165
rect 59 -2199 75 -2182
rect -75 -2215 75 -2199
rect 183 -2199 199 -2182
rect 317 -2182 358 -2165
rect 317 -2199 333 -2182
rect 183 -2215 333 -2199
rect -333 -2273 -183 -2257
rect -333 -2290 -317 -2273
rect -358 -2307 -317 -2290
rect -199 -2290 -183 -2273
rect -75 -2273 75 -2257
rect -75 -2290 -59 -2273
rect -199 -2307 -158 -2290
rect -358 -2354 -158 -2307
rect -100 -2307 -59 -2290
rect 59 -2290 75 -2273
rect 183 -2273 333 -2257
rect 183 -2290 199 -2273
rect 59 -2307 100 -2290
rect -100 -2354 100 -2307
rect 158 -2307 199 -2290
rect 317 -2290 333 -2273
rect 317 -2307 358 -2290
rect 158 -2354 358 -2307
rect -358 -4401 -158 -4354
rect -358 -4418 -317 -4401
rect -333 -4435 -317 -4418
rect -199 -4418 -158 -4401
rect -100 -4401 100 -4354
rect -100 -4418 -59 -4401
rect -199 -4435 -183 -4418
rect -333 -4451 -183 -4435
rect -75 -4435 -59 -4418
rect 59 -4418 100 -4401
rect 158 -4401 358 -4354
rect 158 -4418 199 -4401
rect 59 -4435 75 -4418
rect -75 -4451 75 -4435
rect 183 -4435 199 -4418
rect 317 -4418 358 -4401
rect 317 -4435 333 -4418
rect 183 -4451 333 -4435
<< polycont >>
rect -317 4401 -199 4435
rect -59 4401 59 4435
rect 199 4401 317 4435
rect -317 2273 -199 2307
rect -59 2273 59 2307
rect 199 2273 317 2307
rect -317 2165 -199 2199
rect -59 2165 59 2199
rect 199 2165 317 2199
rect -317 37 -199 71
rect -59 37 59 71
rect 199 37 317 71
rect -317 -71 -199 -37
rect -59 -71 59 -37
rect 199 -71 317 -37
rect -317 -2199 -199 -2165
rect -59 -2199 59 -2165
rect 199 -2199 317 -2165
rect -317 -2307 -199 -2273
rect -59 -2307 59 -2273
rect 199 -2307 317 -2273
rect -317 -4435 -199 -4401
rect -59 -4435 59 -4401
rect 199 -4435 317 -4401
<< locali >>
rect -518 4503 -339 4537
rect 339 4503 518 4537
rect -518 3152 -484 4503
rect -404 4046 -370 4062
rect -404 2646 -370 2662
rect -146 4046 -112 4062
rect -146 2646 -112 2662
rect 112 4046 146 4062
rect 112 2646 146 2662
rect 370 4046 404 4062
rect 370 2646 404 2662
rect 484 3152 518 4503
rect -404 1810 -370 1826
rect -404 410 -370 426
rect -146 1810 -112 1826
rect -146 410 -112 426
rect 112 1810 146 1826
rect 112 410 146 426
rect 370 1810 404 1826
rect 370 410 404 426
rect -404 -426 -370 -410
rect -404 -1826 -370 -1810
rect -146 -426 -112 -410
rect -146 -1826 -112 -1810
rect 112 -426 146 -410
rect 112 -1826 146 -1810
rect 370 -426 404 -410
rect 370 -1826 404 -1810
rect -518 -4503 -484 -3152
rect -404 -2662 -370 -2646
rect -404 -4062 -370 -4046
rect -146 -2662 -112 -2646
rect -146 -4062 -112 -4046
rect 112 -2662 146 -2646
rect 112 -4062 146 -4046
rect 370 -2662 404 -2646
rect 370 -4062 404 -4046
rect 484 -4503 518 -3152
rect -518 -4537 -339 -4503
rect 339 -4537 518 -4503
<< viali >>
rect -339 4503 -295 4537
rect -295 4503 295 4537
rect 295 4503 339 4537
rect -342 4401 -317 4435
rect -317 4401 -199 4435
rect -199 4401 -174 4435
rect -84 4401 -59 4435
rect -59 4401 59 4435
rect 59 4401 84 4435
rect 174 4401 199 4435
rect 199 4401 317 4435
rect 317 4401 342 4435
rect -518 3109 -484 3152
rect -518 -3109 -484 3109
rect -404 2662 -370 4046
rect -146 2662 -112 4046
rect 112 2662 146 4046
rect 370 2662 404 4046
rect 484 3109 518 3152
rect -342 2273 -317 2307
rect -317 2273 -199 2307
rect -199 2273 -174 2307
rect -84 2273 -59 2307
rect -59 2273 59 2307
rect 59 2273 84 2307
rect 174 2273 199 2307
rect 199 2273 317 2307
rect 317 2273 342 2307
rect -342 2165 -317 2199
rect -317 2165 -199 2199
rect -199 2165 -174 2199
rect -84 2165 -59 2199
rect -59 2165 59 2199
rect 59 2165 84 2199
rect 174 2165 199 2199
rect 199 2165 317 2199
rect 317 2165 342 2199
rect -404 426 -370 1810
rect -146 426 -112 1810
rect 112 426 146 1810
rect 370 426 404 1810
rect -342 37 -317 71
rect -317 37 -199 71
rect -199 37 -174 71
rect -84 37 -59 71
rect -59 37 59 71
rect 59 37 84 71
rect 174 37 199 71
rect 199 37 317 71
rect 317 37 342 71
rect -342 -71 -317 -37
rect -317 -71 -199 -37
rect -199 -71 -174 -37
rect -84 -71 -59 -37
rect -59 -71 59 -37
rect 59 -71 84 -37
rect 174 -71 199 -37
rect 199 -71 317 -37
rect 317 -71 342 -37
rect -404 -1810 -370 -426
rect -146 -1810 -112 -426
rect 112 -1810 146 -426
rect 370 -1810 404 -426
rect -342 -2199 -317 -2165
rect -317 -2199 -199 -2165
rect -199 -2199 -174 -2165
rect -84 -2199 -59 -2165
rect -59 -2199 59 -2165
rect 59 -2199 84 -2165
rect 174 -2199 199 -2165
rect 199 -2199 317 -2165
rect 317 -2199 342 -2165
rect -342 -2307 -317 -2273
rect -317 -2307 -199 -2273
rect -199 -2307 -174 -2273
rect -84 -2307 -59 -2273
rect -59 -2307 59 -2273
rect 59 -2307 84 -2273
rect 174 -2307 199 -2273
rect 199 -2307 317 -2273
rect 317 -2307 342 -2273
rect -518 -3152 -484 -3109
rect -404 -4046 -370 -2662
rect -146 -4046 -112 -2662
rect 112 -4046 146 -2662
rect 370 -4046 404 -2662
rect 484 -3109 518 3109
rect 484 -3152 518 -3109
rect -342 -4435 -317 -4401
rect -317 -4435 -199 -4401
rect -199 -4435 -174 -4401
rect -84 -4435 -59 -4401
rect -59 -4435 59 -4401
rect 59 -4435 84 -4401
rect 174 -4435 199 -4401
rect 199 -4435 317 -4401
rect 317 -4435 342 -4401
rect -339 -4537 -295 -4503
rect -295 -4537 295 -4503
rect 295 -4537 339 -4503
<< metal1 >>
rect -351 4537 351 4543
rect -351 4503 -339 4537
rect 339 4503 351 4537
rect -351 4497 351 4503
rect -354 4435 -162 4441
rect -354 4401 -342 4435
rect -174 4401 -162 4435
rect -354 4395 -162 4401
rect -96 4435 96 4441
rect -96 4401 -84 4435
rect 84 4401 96 4435
rect -96 4395 96 4401
rect 162 4435 354 4441
rect 162 4401 174 4435
rect 342 4401 354 4435
rect 162 4395 354 4401
rect -410 4046 -364 4058
rect -524 3152 -478 3164
rect -524 -3152 -518 3152
rect -484 -3152 -478 3152
rect -410 2662 -404 4046
rect -370 2662 -364 4046
rect -410 2650 -364 2662
rect -152 4046 -106 4058
rect -152 2662 -146 4046
rect -112 2662 -106 4046
rect -152 2650 -106 2662
rect 106 4046 152 4058
rect 106 2662 112 4046
rect 146 2662 152 4046
rect 106 2650 152 2662
rect 364 4046 410 4058
rect 364 2662 370 4046
rect 404 2662 410 4046
rect 364 2650 410 2662
rect 478 3152 524 3164
rect -354 2307 -162 2313
rect -354 2273 -342 2307
rect -174 2273 -162 2307
rect -354 2267 -162 2273
rect -96 2307 96 2313
rect -96 2273 -84 2307
rect 84 2273 96 2307
rect -96 2267 96 2273
rect 162 2307 354 2313
rect 162 2273 174 2307
rect 342 2273 354 2307
rect 162 2267 354 2273
rect -354 2199 -162 2205
rect -354 2165 -342 2199
rect -174 2165 -162 2199
rect -354 2159 -162 2165
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect 162 2199 354 2205
rect 162 2165 174 2199
rect 342 2165 354 2199
rect 162 2159 354 2165
rect -410 1810 -364 1822
rect -410 426 -404 1810
rect -370 426 -364 1810
rect -410 414 -364 426
rect -152 1810 -106 1822
rect -152 426 -146 1810
rect -112 426 -106 1810
rect -152 414 -106 426
rect 106 1810 152 1822
rect 106 426 112 1810
rect 146 426 152 1810
rect 106 414 152 426
rect 364 1810 410 1822
rect 364 426 370 1810
rect 404 426 410 1810
rect 364 414 410 426
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect -410 -426 -364 -414
rect -410 -1810 -404 -426
rect -370 -1810 -364 -426
rect -410 -1822 -364 -1810
rect -152 -426 -106 -414
rect -152 -1810 -146 -426
rect -112 -1810 -106 -426
rect -152 -1822 -106 -1810
rect 106 -426 152 -414
rect 106 -1810 112 -426
rect 146 -1810 152 -426
rect 106 -1822 152 -1810
rect 364 -426 410 -414
rect 364 -1810 370 -426
rect 404 -1810 410 -426
rect 364 -1822 410 -1810
rect -354 -2165 -162 -2159
rect -354 -2199 -342 -2165
rect -174 -2199 -162 -2165
rect -354 -2205 -162 -2199
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
rect 162 -2165 354 -2159
rect 162 -2199 174 -2165
rect 342 -2199 354 -2165
rect 162 -2205 354 -2199
rect -354 -2273 -162 -2267
rect -354 -2307 -342 -2273
rect -174 -2307 -162 -2273
rect -354 -2313 -162 -2307
rect -96 -2273 96 -2267
rect -96 -2307 -84 -2273
rect 84 -2307 96 -2273
rect -96 -2313 96 -2307
rect 162 -2273 354 -2267
rect 162 -2307 174 -2273
rect 342 -2307 354 -2273
rect 162 -2313 354 -2307
rect -524 -3164 -478 -3152
rect -410 -2662 -364 -2650
rect -410 -4046 -404 -2662
rect -370 -4046 -364 -2662
rect -410 -4058 -364 -4046
rect -152 -2662 -106 -2650
rect -152 -4046 -146 -2662
rect -112 -4046 -106 -2662
rect -152 -4058 -106 -4046
rect 106 -2662 152 -2650
rect 106 -4046 112 -2662
rect 146 -4046 152 -2662
rect 106 -4058 152 -4046
rect 364 -2662 410 -2650
rect 364 -4046 370 -2662
rect 404 -4046 410 -2662
rect 478 -3152 484 3152
rect 518 -3152 524 3152
rect 478 -3164 524 -3152
rect 364 -4058 410 -4046
rect -354 -4401 -162 -4395
rect -354 -4435 -342 -4401
rect -174 -4435 -162 -4401
rect -354 -4441 -162 -4435
rect -96 -4401 96 -4395
rect -96 -4435 -84 -4401
rect 84 -4435 96 -4401
rect -96 -4441 96 -4435
rect 162 -4401 354 -4395
rect 162 -4435 174 -4401
rect 342 -4435 354 -4401
rect 162 -4441 354 -4435
rect -351 -4503 351 -4497
rect -351 -4537 -339 -4503
rect 339 -4537 351 -4503
rect -351 -4543 351 -4537
<< properties >>
string FIXED_BBOX -501 -4520 501 4520
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 4 nf 3 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
