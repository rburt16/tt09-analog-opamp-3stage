magic
tech sky130A
magscale 1 2
timestamp 1730563144
<< nwell >>
rect -554 -2337 554 2337
<< pmos >>
rect -358 118 -158 2118
rect -100 118 100 2118
rect 158 118 358 2118
rect -358 -2118 -158 -118
rect -100 -2118 100 -118
rect 158 -2118 358 -118
<< pdiff >>
rect -416 1810 -358 2118
rect -416 426 -404 1810
rect -370 426 -358 1810
rect -416 118 -358 426
rect -158 1810 -100 2118
rect -158 426 -146 1810
rect -112 426 -100 1810
rect -158 118 -100 426
rect 100 1810 158 2118
rect 100 426 112 1810
rect 146 426 158 1810
rect 100 118 158 426
rect 358 1810 416 2118
rect 358 426 370 1810
rect 404 426 416 1810
rect 358 118 416 426
rect -416 -426 -358 -118
rect -416 -1810 -404 -426
rect -370 -1810 -358 -426
rect -416 -2118 -358 -1810
rect -158 -426 -100 -118
rect -158 -1810 -146 -426
rect -112 -1810 -100 -426
rect -158 -2118 -100 -1810
rect 100 -426 158 -118
rect 100 -1810 112 -426
rect 146 -1810 158 -426
rect 100 -2118 158 -1810
rect 358 -426 416 -118
rect 358 -1810 370 -426
rect 404 -1810 416 -426
rect 358 -2118 416 -1810
<< pdiffc >>
rect -404 426 -370 1810
rect -146 426 -112 1810
rect 112 426 146 1810
rect 370 426 404 1810
rect -404 -1810 -370 -426
rect -146 -1810 -112 -426
rect 112 -1810 146 -426
rect 370 -1810 404 -426
<< nsubdiff >>
rect -518 2267 -295 2301
rect 295 2267 518 2301
rect -518 1544 -484 2267
rect 484 1544 518 2267
rect -518 -2267 -484 -1544
rect 484 -2267 518 -1544
rect -518 -2301 -295 -2267
rect 295 -2301 518 -2267
<< nsubdiffcont >>
rect -295 2267 295 2301
rect -518 -1544 -484 1544
rect 484 -1544 518 1544
rect -295 -2301 295 -2267
<< poly >>
rect -333 2199 -183 2215
rect -333 2182 -317 2199
rect -358 2165 -317 2182
rect -199 2182 -183 2199
rect -75 2199 75 2215
rect -75 2182 -59 2199
rect -199 2165 -158 2182
rect -358 2118 -158 2165
rect -100 2165 -59 2182
rect 59 2182 75 2199
rect 183 2199 333 2215
rect 183 2182 199 2199
rect 59 2165 100 2182
rect -100 2118 100 2165
rect 158 2165 199 2182
rect 317 2182 333 2199
rect 317 2165 358 2182
rect 158 2118 358 2165
rect -358 71 -158 118
rect -358 54 -317 71
rect -333 37 -317 54
rect -199 54 -158 71
rect -100 71 100 118
rect -100 54 -59 71
rect -199 37 -183 54
rect -333 21 -183 37
rect -75 37 -59 54
rect 59 54 100 71
rect 158 71 358 118
rect 158 54 199 71
rect 59 37 75 54
rect -75 21 75 37
rect 183 37 199 54
rect 317 54 358 71
rect 317 37 333 54
rect 183 21 333 37
rect -333 -37 -183 -21
rect -333 -54 -317 -37
rect -358 -71 -317 -54
rect -199 -54 -183 -37
rect -75 -37 75 -21
rect -75 -54 -59 -37
rect -199 -71 -158 -54
rect -358 -118 -158 -71
rect -100 -71 -59 -54
rect 59 -54 75 -37
rect 183 -37 333 -21
rect 183 -54 199 -37
rect 59 -71 100 -54
rect -100 -118 100 -71
rect 158 -71 199 -54
rect 317 -54 333 -37
rect 317 -71 358 -54
rect 158 -118 358 -71
rect -358 -2165 -158 -2118
rect -358 -2182 -317 -2165
rect -333 -2199 -317 -2182
rect -199 -2182 -158 -2165
rect -100 -2165 100 -2118
rect -100 -2182 -59 -2165
rect -199 -2199 -183 -2182
rect -333 -2215 -183 -2199
rect -75 -2199 -59 -2182
rect 59 -2182 100 -2165
rect 158 -2165 358 -2118
rect 158 -2182 199 -2165
rect 59 -2199 75 -2182
rect -75 -2215 75 -2199
rect 183 -2199 199 -2182
rect 317 -2182 358 -2165
rect 317 -2199 333 -2182
rect 183 -2215 333 -2199
<< polycont >>
rect -317 2165 -199 2199
rect -59 2165 59 2199
rect 199 2165 317 2199
rect -317 37 -199 71
rect -59 37 59 71
rect 199 37 317 71
rect -317 -71 -199 -37
rect -59 -71 59 -37
rect 199 -71 317 -37
rect -317 -2199 -199 -2165
rect -59 -2199 59 -2165
rect 199 -2199 317 -2165
<< locali >>
rect -518 2267 -339 2301
rect 339 2267 518 2301
rect -518 1587 -484 2267
rect -404 1810 -370 1826
rect -404 410 -370 426
rect -146 1810 -112 1826
rect -146 410 -112 426
rect 112 1810 146 1826
rect 112 410 146 426
rect 370 1810 404 1826
rect 370 410 404 426
rect 484 1587 518 2267
rect -518 -2267 -484 -1587
rect -404 -426 -370 -410
rect -404 -1826 -370 -1810
rect -146 -426 -112 -410
rect -146 -1826 -112 -1810
rect 112 -426 146 -410
rect 112 -1826 146 -1810
rect 370 -426 404 -410
rect 370 -1826 404 -1810
rect 484 -2267 518 -1587
rect -518 -2301 -339 -2267
rect 339 -2301 518 -2267
<< viali >>
rect -339 2267 -295 2301
rect -295 2267 295 2301
rect 295 2267 339 2301
rect -342 2165 -317 2199
rect -317 2165 -199 2199
rect -199 2165 -174 2199
rect -84 2165 -59 2199
rect -59 2165 59 2199
rect 59 2165 84 2199
rect 174 2165 199 2199
rect 199 2165 317 2199
rect 317 2165 342 2199
rect -518 1544 -484 1587
rect -518 -1544 -484 1544
rect -404 426 -370 1810
rect -146 426 -112 1810
rect 112 426 146 1810
rect 370 426 404 1810
rect 484 1544 518 1587
rect -342 37 -317 71
rect -317 37 -199 71
rect -199 37 -174 71
rect -84 37 -59 71
rect -59 37 59 71
rect 59 37 84 71
rect 174 37 199 71
rect 199 37 317 71
rect 317 37 342 71
rect -342 -71 -317 -37
rect -317 -71 -199 -37
rect -199 -71 -174 -37
rect -84 -71 -59 -37
rect -59 -71 59 -37
rect 59 -71 84 -37
rect 174 -71 199 -37
rect 199 -71 317 -37
rect 317 -71 342 -37
rect -518 -1587 -484 -1544
rect -404 -1810 -370 -426
rect -146 -1810 -112 -426
rect 112 -1810 146 -426
rect 370 -1810 404 -426
rect 484 -1544 518 1544
rect 484 -1587 518 -1544
rect -342 -2199 -317 -2165
rect -317 -2199 -199 -2165
rect -199 -2199 -174 -2165
rect -84 -2199 -59 -2165
rect -59 -2199 59 -2165
rect 59 -2199 84 -2165
rect 174 -2199 199 -2165
rect 199 -2199 317 -2165
rect 317 -2199 342 -2165
rect -339 -2301 -295 -2267
rect -295 -2301 295 -2267
rect 295 -2301 339 -2267
<< metal1 >>
rect -351 2301 351 2307
rect -351 2267 -339 2301
rect 339 2267 351 2301
rect -351 2261 351 2267
rect -354 2199 -162 2205
rect -354 2165 -342 2199
rect -174 2165 -162 2199
rect -354 2159 -162 2165
rect -96 2199 96 2205
rect -96 2165 -84 2199
rect 84 2165 96 2199
rect -96 2159 96 2165
rect 162 2199 354 2205
rect 162 2165 174 2199
rect 342 2165 354 2199
rect 162 2159 354 2165
rect -410 1810 -364 1822
rect -524 1587 -478 1599
rect -524 -1587 -518 1587
rect -484 -1587 -478 1587
rect -410 426 -404 1810
rect -370 426 -364 1810
rect -410 414 -364 426
rect -152 1810 -106 1822
rect -152 426 -146 1810
rect -112 426 -106 1810
rect -152 414 -106 426
rect 106 1810 152 1822
rect 106 426 112 1810
rect 146 426 152 1810
rect 106 414 152 426
rect 364 1810 410 1822
rect 364 426 370 1810
rect 404 426 410 1810
rect 364 414 410 426
rect 478 1587 524 1599
rect -354 71 -162 77
rect -354 37 -342 71
rect -174 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 174 71
rect 342 37 354 71
rect 162 31 354 37
rect -354 -37 -162 -31
rect -354 -71 -342 -37
rect -174 -71 -162 -37
rect -354 -77 -162 -71
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect 162 -37 354 -31
rect 162 -71 174 -37
rect 342 -71 354 -37
rect 162 -77 354 -71
rect -524 -1599 -478 -1587
rect -410 -426 -364 -414
rect -410 -1810 -404 -426
rect -370 -1810 -364 -426
rect -410 -1822 -364 -1810
rect -152 -426 -106 -414
rect -152 -1810 -146 -426
rect -112 -1810 -106 -426
rect -152 -1822 -106 -1810
rect 106 -426 152 -414
rect 106 -1810 112 -426
rect 146 -1810 152 -426
rect 106 -1822 152 -1810
rect 364 -426 410 -414
rect 364 -1810 370 -426
rect 404 -1810 410 -426
rect 478 -1587 484 1587
rect 518 -1587 524 1587
rect 478 -1599 524 -1587
rect 364 -1822 410 -1810
rect -354 -2165 -162 -2159
rect -354 -2199 -342 -2165
rect -174 -2199 -162 -2165
rect -354 -2205 -162 -2199
rect -96 -2165 96 -2159
rect -96 -2199 -84 -2165
rect 84 -2199 96 -2165
rect -96 -2205 96 -2199
rect 162 -2165 354 -2159
rect 162 -2199 174 -2165
rect 342 -2199 354 -2165
rect 162 -2205 354 -2199
rect -351 -2267 351 -2261
rect -351 -2301 -339 -2267
rect 339 -2301 351 -2267
rect -351 -2307 351 -2301
<< properties >>
string FIXED_BBOX -501 -2284 501 2284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 2 nf 3 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
