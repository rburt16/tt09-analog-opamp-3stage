magic
tech sky130A
magscale 1 2
timestamp 1730569394
<< error_p >>
rect -1055 681 -993 687
rect -927 681 -865 687
rect -799 681 -737 687
rect -671 681 -609 687
rect -543 681 -481 687
rect -415 681 -353 687
rect -287 681 -225 687
rect -159 681 -97 687
rect -31 681 31 687
rect 97 681 159 687
rect 225 681 287 687
rect 353 681 415 687
rect 481 681 543 687
rect 609 681 671 687
rect 737 681 799 687
rect 865 681 927 687
rect 993 681 1055 687
rect -1055 647 -1043 681
rect -927 647 -915 681
rect -799 647 -787 681
rect -671 647 -659 681
rect -543 647 -531 681
rect -415 647 -403 681
rect -287 647 -275 681
rect -159 647 -147 681
rect -31 647 -19 681
rect 97 647 109 681
rect 225 647 237 681
rect 353 647 365 681
rect 481 647 493 681
rect 609 647 621 681
rect 737 647 749 681
rect 865 647 877 681
rect 993 647 1005 681
rect -1055 641 -993 647
rect -927 641 -865 647
rect -799 641 -737 647
rect -671 641 -609 647
rect -543 641 -481 647
rect -415 641 -353 647
rect -287 641 -225 647
rect -159 641 -97 647
rect -31 641 31 647
rect 97 641 159 647
rect 225 641 287 647
rect 353 641 415 647
rect 481 641 543 647
rect 609 641 671 647
rect 737 641 799 647
rect 865 641 927 647
rect 993 641 1055 647
rect -1055 71 -993 77
rect -927 71 -865 77
rect -799 71 -737 77
rect -671 71 -609 77
rect -543 71 -481 77
rect -415 71 -353 77
rect -287 71 -225 77
rect -159 71 -97 77
rect -31 71 31 77
rect 97 71 159 77
rect 225 71 287 77
rect 353 71 415 77
rect 481 71 543 77
rect 609 71 671 77
rect 737 71 799 77
rect 865 71 927 77
rect 993 71 1055 77
rect -1055 37 -1043 71
rect -927 37 -915 71
rect -799 37 -787 71
rect -671 37 -659 71
rect -543 37 -531 71
rect -415 37 -403 71
rect -287 37 -275 71
rect -159 37 -147 71
rect -31 37 -19 71
rect 97 37 109 71
rect 225 37 237 71
rect 353 37 365 71
rect 481 37 493 71
rect 609 37 621 71
rect 737 37 749 71
rect 865 37 877 71
rect 993 37 1005 71
rect -1055 31 -993 37
rect -927 31 -865 37
rect -799 31 -737 37
rect -671 31 -609 37
rect -543 31 -481 37
rect -415 31 -353 37
rect -287 31 -225 37
rect -159 31 -97 37
rect -31 31 31 37
rect 97 31 159 37
rect 225 31 287 37
rect 353 31 415 37
rect 481 31 543 37
rect 609 31 671 37
rect 737 31 799 37
rect 865 31 927 37
rect 993 31 1055 37
rect -1055 -37 -993 -31
rect -927 -37 -865 -31
rect -799 -37 -737 -31
rect -671 -37 -609 -31
rect -543 -37 -481 -31
rect -415 -37 -353 -31
rect -287 -37 -225 -31
rect -159 -37 -97 -31
rect -31 -37 31 -31
rect 97 -37 159 -31
rect 225 -37 287 -31
rect 353 -37 415 -31
rect 481 -37 543 -31
rect 609 -37 671 -31
rect 737 -37 799 -31
rect 865 -37 927 -31
rect 993 -37 1055 -31
rect -1055 -71 -1043 -37
rect -927 -71 -915 -37
rect -799 -71 -787 -37
rect -671 -71 -659 -37
rect -543 -71 -531 -37
rect -415 -71 -403 -37
rect -287 -71 -275 -37
rect -159 -71 -147 -37
rect -31 -71 -19 -37
rect 97 -71 109 -37
rect 225 -71 237 -37
rect 353 -71 365 -37
rect 481 -71 493 -37
rect 609 -71 621 -37
rect 737 -71 749 -37
rect 865 -71 877 -37
rect 993 -71 1005 -37
rect -1055 -77 -993 -71
rect -927 -77 -865 -71
rect -799 -77 -737 -71
rect -671 -77 -609 -71
rect -543 -77 -481 -71
rect -415 -77 -353 -71
rect -287 -77 -225 -71
rect -159 -77 -97 -71
rect -31 -77 31 -71
rect 97 -77 159 -71
rect 225 -77 287 -71
rect 353 -77 415 -71
rect 481 -77 543 -71
rect 609 -77 671 -71
rect 737 -77 799 -71
rect 865 -77 927 -71
rect 993 -77 1055 -71
rect -1055 -647 -993 -641
rect -927 -647 -865 -641
rect -799 -647 -737 -641
rect -671 -647 -609 -641
rect -543 -647 -481 -641
rect -415 -647 -353 -641
rect -287 -647 -225 -641
rect -159 -647 -97 -641
rect -31 -647 31 -641
rect 97 -647 159 -641
rect 225 -647 287 -641
rect 353 -647 415 -641
rect 481 -647 543 -641
rect 609 -647 671 -641
rect 737 -647 799 -641
rect 865 -647 927 -641
rect 993 -647 1055 -641
rect -1055 -681 -1043 -647
rect -927 -681 -915 -647
rect -799 -681 -787 -647
rect -671 -681 -659 -647
rect -543 -681 -531 -647
rect -415 -681 -403 -647
rect -287 -681 -275 -647
rect -159 -681 -147 -647
rect -31 -681 -19 -647
rect 97 -681 109 -647
rect 225 -681 237 -647
rect 353 -681 365 -647
rect 481 -681 493 -647
rect 609 -681 621 -647
rect 737 -681 749 -647
rect 865 -681 877 -647
rect 993 -681 1005 -647
rect -1055 -687 -993 -681
rect -927 -687 -865 -681
rect -799 -687 -737 -681
rect -671 -687 -609 -681
rect -543 -687 -481 -681
rect -415 -687 -353 -681
rect -287 -687 -225 -681
rect -159 -687 -97 -681
rect -31 -687 31 -681
rect 97 -687 159 -681
rect 225 -687 287 -681
rect 353 -687 415 -681
rect 481 -687 543 -681
rect 609 -687 671 -681
rect 737 -687 799 -681
rect 865 -687 927 -681
rect 993 -687 1055 -681
<< pwell >>
rect -1255 -819 1255 819
<< nmoslvt >>
rect -1059 109 -989 609
rect -931 109 -861 609
rect -803 109 -733 609
rect -675 109 -605 609
rect -547 109 -477 609
rect -419 109 -349 609
rect -291 109 -221 609
rect -163 109 -93 609
rect -35 109 35 609
rect 93 109 163 609
rect 221 109 291 609
rect 349 109 419 609
rect 477 109 547 609
rect 605 109 675 609
rect 733 109 803 609
rect 861 109 931 609
rect 989 109 1059 609
rect -1059 -609 -989 -109
rect -931 -609 -861 -109
rect -803 -609 -733 -109
rect -675 -609 -605 -109
rect -547 -609 -477 -109
rect -419 -609 -349 -109
rect -291 -609 -221 -109
rect -163 -609 -93 -109
rect -35 -609 35 -109
rect 93 -609 163 -109
rect 221 -609 291 -109
rect 349 -609 419 -109
rect 477 -609 547 -109
rect 605 -609 675 -109
rect 733 -609 803 -109
rect 861 -609 931 -109
rect 989 -609 1059 -109
<< ndiff >>
rect -1117 407 -1059 609
rect -1117 311 -1105 407
rect -1071 311 -1059 407
rect -1117 109 -1059 311
rect -989 407 -931 609
rect -989 311 -977 407
rect -943 311 -931 407
rect -989 109 -931 311
rect -861 407 -803 609
rect -861 311 -849 407
rect -815 311 -803 407
rect -861 109 -803 311
rect -733 407 -675 609
rect -733 311 -721 407
rect -687 311 -675 407
rect -733 109 -675 311
rect -605 407 -547 609
rect -605 311 -593 407
rect -559 311 -547 407
rect -605 109 -547 311
rect -477 407 -419 609
rect -477 311 -465 407
rect -431 311 -419 407
rect -477 109 -419 311
rect -349 407 -291 609
rect -349 311 -337 407
rect -303 311 -291 407
rect -349 109 -291 311
rect -221 407 -163 609
rect -221 311 -209 407
rect -175 311 -163 407
rect -221 109 -163 311
rect -93 407 -35 609
rect -93 311 -81 407
rect -47 311 -35 407
rect -93 109 -35 311
rect 35 407 93 609
rect 35 311 47 407
rect 81 311 93 407
rect 35 109 93 311
rect 163 407 221 609
rect 163 311 175 407
rect 209 311 221 407
rect 163 109 221 311
rect 291 407 349 609
rect 291 311 303 407
rect 337 311 349 407
rect 291 109 349 311
rect 419 407 477 609
rect 419 311 431 407
rect 465 311 477 407
rect 419 109 477 311
rect 547 407 605 609
rect 547 311 559 407
rect 593 311 605 407
rect 547 109 605 311
rect 675 407 733 609
rect 675 311 687 407
rect 721 311 733 407
rect 675 109 733 311
rect 803 407 861 609
rect 803 311 815 407
rect 849 311 861 407
rect 803 109 861 311
rect 931 407 989 609
rect 931 311 943 407
rect 977 311 989 407
rect 931 109 989 311
rect 1059 407 1117 609
rect 1059 311 1071 407
rect 1105 311 1117 407
rect 1059 109 1117 311
rect -1117 -311 -1059 -109
rect -1117 -407 -1105 -311
rect -1071 -407 -1059 -311
rect -1117 -609 -1059 -407
rect -989 -311 -931 -109
rect -989 -407 -977 -311
rect -943 -407 -931 -311
rect -989 -609 -931 -407
rect -861 -311 -803 -109
rect -861 -407 -849 -311
rect -815 -407 -803 -311
rect -861 -609 -803 -407
rect -733 -311 -675 -109
rect -733 -407 -721 -311
rect -687 -407 -675 -311
rect -733 -609 -675 -407
rect -605 -311 -547 -109
rect -605 -407 -593 -311
rect -559 -407 -547 -311
rect -605 -609 -547 -407
rect -477 -311 -419 -109
rect -477 -407 -465 -311
rect -431 -407 -419 -311
rect -477 -609 -419 -407
rect -349 -311 -291 -109
rect -349 -407 -337 -311
rect -303 -407 -291 -311
rect -349 -609 -291 -407
rect -221 -311 -163 -109
rect -221 -407 -209 -311
rect -175 -407 -163 -311
rect -221 -609 -163 -407
rect -93 -311 -35 -109
rect -93 -407 -81 -311
rect -47 -407 -35 -311
rect -93 -609 -35 -407
rect 35 -311 93 -109
rect 35 -407 47 -311
rect 81 -407 93 -311
rect 35 -609 93 -407
rect 163 -311 221 -109
rect 163 -407 175 -311
rect 209 -407 221 -311
rect 163 -609 221 -407
rect 291 -311 349 -109
rect 291 -407 303 -311
rect 337 -407 349 -311
rect 291 -609 349 -407
rect 419 -311 477 -109
rect 419 -407 431 -311
rect 465 -407 477 -311
rect 419 -609 477 -407
rect 547 -311 605 -109
rect 547 -407 559 -311
rect 593 -407 605 -311
rect 547 -609 605 -407
rect 675 -311 733 -109
rect 675 -407 687 -311
rect 721 -407 733 -311
rect 675 -609 733 -407
rect 803 -311 861 -109
rect 803 -407 815 -311
rect 849 -407 861 -311
rect 803 -609 861 -407
rect 931 -311 989 -109
rect 931 -407 943 -311
rect 977 -407 989 -311
rect 931 -609 989 -407
rect 1059 -311 1117 -109
rect 1059 -407 1071 -311
rect 1105 -407 1117 -311
rect 1059 -609 1117 -407
<< ndiffc >>
rect -1105 311 -1071 407
rect -977 311 -943 407
rect -849 311 -815 407
rect -721 311 -687 407
rect -593 311 -559 407
rect -465 311 -431 407
rect -337 311 -303 407
rect -209 311 -175 407
rect -81 311 -47 407
rect 47 311 81 407
rect 175 311 209 407
rect 303 311 337 407
rect 431 311 465 407
rect 559 311 593 407
rect 687 311 721 407
rect 815 311 849 407
rect 943 311 977 407
rect 1071 311 1105 407
rect -1105 -407 -1071 -311
rect -977 -407 -943 -311
rect -849 -407 -815 -311
rect -721 -407 -687 -311
rect -593 -407 -559 -311
rect -465 -407 -431 -311
rect -337 -407 -303 -311
rect -209 -407 -175 -311
rect -81 -407 -47 -311
rect 47 -407 81 -311
rect 175 -407 209 -311
rect 303 -407 337 -311
rect 431 -407 465 -311
rect 559 -407 593 -311
rect 687 -407 721 -311
rect 815 -407 849 -311
rect 943 -407 977 -311
rect 1071 -407 1105 -311
<< psubdiff >>
rect -1219 749 1219 783
rect -1219 481 -1185 749
rect -1219 -749 -1185 -481
rect 1185 -749 1219 749
rect -1219 -783 1219 -749
<< psubdiffcont >>
rect -1219 -481 -1185 481
<< poly >>
rect -1057 681 -991 697
rect -1057 664 -1041 681
rect -1059 647 -1041 664
rect -1007 664 -991 681
rect -929 681 -863 697
rect -929 664 -913 681
rect -1007 647 -989 664
rect -1059 609 -989 647
rect -931 647 -913 664
rect -879 664 -863 681
rect -801 681 -735 697
rect -801 664 -785 681
rect -879 647 -861 664
rect -931 609 -861 647
rect -803 647 -785 664
rect -751 664 -735 681
rect -673 681 -607 697
rect -673 664 -657 681
rect -751 647 -733 664
rect -803 609 -733 647
rect -675 647 -657 664
rect -623 664 -607 681
rect -545 681 -479 697
rect -545 664 -529 681
rect -623 647 -605 664
rect -675 609 -605 647
rect -547 647 -529 664
rect -495 664 -479 681
rect -417 681 -351 697
rect -417 664 -401 681
rect -495 647 -477 664
rect -547 609 -477 647
rect -419 647 -401 664
rect -367 664 -351 681
rect -289 681 -223 697
rect -289 664 -273 681
rect -367 647 -349 664
rect -419 609 -349 647
rect -291 647 -273 664
rect -239 664 -223 681
rect -161 681 -95 697
rect -161 664 -145 681
rect -239 647 -221 664
rect -291 609 -221 647
rect -163 647 -145 664
rect -111 664 -95 681
rect -33 681 33 697
rect -33 664 -17 681
rect -111 647 -93 664
rect -163 609 -93 647
rect -35 647 -17 664
rect 17 664 33 681
rect 95 681 161 697
rect 95 664 111 681
rect 17 647 35 664
rect -35 609 35 647
rect 93 647 111 664
rect 145 664 161 681
rect 223 681 289 697
rect 223 664 239 681
rect 145 647 163 664
rect 93 609 163 647
rect 221 647 239 664
rect 273 664 289 681
rect 351 681 417 697
rect 351 664 367 681
rect 273 647 291 664
rect 221 609 291 647
rect 349 647 367 664
rect 401 664 417 681
rect 479 681 545 697
rect 479 664 495 681
rect 401 647 419 664
rect 349 609 419 647
rect 477 647 495 664
rect 529 664 545 681
rect 607 681 673 697
rect 607 664 623 681
rect 529 647 547 664
rect 477 609 547 647
rect 605 647 623 664
rect 657 664 673 681
rect 735 681 801 697
rect 735 664 751 681
rect 657 647 675 664
rect 605 609 675 647
rect 733 647 751 664
rect 785 664 801 681
rect 863 681 929 697
rect 863 664 879 681
rect 785 647 803 664
rect 733 609 803 647
rect 861 647 879 664
rect 913 664 929 681
rect 991 681 1057 697
rect 991 664 1007 681
rect 913 647 931 664
rect 861 609 931 647
rect 989 647 1007 664
rect 1041 664 1057 681
rect 1041 647 1059 664
rect 989 609 1059 647
rect -1059 71 -989 109
rect -1059 54 -1041 71
rect -1057 37 -1041 54
rect -1007 54 -989 71
rect -931 71 -861 109
rect -931 54 -913 71
rect -1007 37 -991 54
rect -1057 21 -991 37
rect -929 37 -913 54
rect -879 54 -861 71
rect -803 71 -733 109
rect -803 54 -785 71
rect -879 37 -863 54
rect -929 21 -863 37
rect -801 37 -785 54
rect -751 54 -733 71
rect -675 71 -605 109
rect -675 54 -657 71
rect -751 37 -735 54
rect -801 21 -735 37
rect -673 37 -657 54
rect -623 54 -605 71
rect -547 71 -477 109
rect -547 54 -529 71
rect -623 37 -607 54
rect -673 21 -607 37
rect -545 37 -529 54
rect -495 54 -477 71
rect -419 71 -349 109
rect -419 54 -401 71
rect -495 37 -479 54
rect -545 21 -479 37
rect -417 37 -401 54
rect -367 54 -349 71
rect -291 71 -221 109
rect -291 54 -273 71
rect -367 37 -351 54
rect -417 21 -351 37
rect -289 37 -273 54
rect -239 54 -221 71
rect -163 71 -93 109
rect -163 54 -145 71
rect -239 37 -223 54
rect -289 21 -223 37
rect -161 37 -145 54
rect -111 54 -93 71
rect -35 71 35 109
rect -35 54 -17 71
rect -111 37 -95 54
rect -161 21 -95 37
rect -33 37 -17 54
rect 17 54 35 71
rect 93 71 163 109
rect 93 54 111 71
rect 17 37 33 54
rect -33 21 33 37
rect 95 37 111 54
rect 145 54 163 71
rect 221 71 291 109
rect 221 54 239 71
rect 145 37 161 54
rect 95 21 161 37
rect 223 37 239 54
rect 273 54 291 71
rect 349 71 419 109
rect 349 54 367 71
rect 273 37 289 54
rect 223 21 289 37
rect 351 37 367 54
rect 401 54 419 71
rect 477 71 547 109
rect 477 54 495 71
rect 401 37 417 54
rect 351 21 417 37
rect 479 37 495 54
rect 529 54 547 71
rect 605 71 675 109
rect 605 54 623 71
rect 529 37 545 54
rect 479 21 545 37
rect 607 37 623 54
rect 657 54 675 71
rect 733 71 803 109
rect 733 54 751 71
rect 657 37 673 54
rect 607 21 673 37
rect 735 37 751 54
rect 785 54 803 71
rect 861 71 931 109
rect 861 54 879 71
rect 785 37 801 54
rect 735 21 801 37
rect 863 37 879 54
rect 913 54 931 71
rect 989 71 1059 109
rect 989 54 1007 71
rect 913 37 929 54
rect 863 21 929 37
rect 991 37 1007 54
rect 1041 54 1059 71
rect 1041 37 1057 54
rect 991 21 1057 37
rect -1057 -37 -991 -21
rect -1057 -54 -1041 -37
rect -1059 -71 -1041 -54
rect -1007 -54 -991 -37
rect -929 -37 -863 -21
rect -929 -54 -913 -37
rect -1007 -71 -989 -54
rect -1059 -109 -989 -71
rect -931 -71 -913 -54
rect -879 -54 -863 -37
rect -801 -37 -735 -21
rect -801 -54 -785 -37
rect -879 -71 -861 -54
rect -931 -109 -861 -71
rect -803 -71 -785 -54
rect -751 -54 -735 -37
rect -673 -37 -607 -21
rect -673 -54 -657 -37
rect -751 -71 -733 -54
rect -803 -109 -733 -71
rect -675 -71 -657 -54
rect -623 -54 -607 -37
rect -545 -37 -479 -21
rect -545 -54 -529 -37
rect -623 -71 -605 -54
rect -675 -109 -605 -71
rect -547 -71 -529 -54
rect -495 -54 -479 -37
rect -417 -37 -351 -21
rect -417 -54 -401 -37
rect -495 -71 -477 -54
rect -547 -109 -477 -71
rect -419 -71 -401 -54
rect -367 -54 -351 -37
rect -289 -37 -223 -21
rect -289 -54 -273 -37
rect -367 -71 -349 -54
rect -419 -109 -349 -71
rect -291 -71 -273 -54
rect -239 -54 -223 -37
rect -161 -37 -95 -21
rect -161 -54 -145 -37
rect -239 -71 -221 -54
rect -291 -109 -221 -71
rect -163 -71 -145 -54
rect -111 -54 -95 -37
rect -33 -37 33 -21
rect -33 -54 -17 -37
rect -111 -71 -93 -54
rect -163 -109 -93 -71
rect -35 -71 -17 -54
rect 17 -54 33 -37
rect 95 -37 161 -21
rect 95 -54 111 -37
rect 17 -71 35 -54
rect -35 -109 35 -71
rect 93 -71 111 -54
rect 145 -54 161 -37
rect 223 -37 289 -21
rect 223 -54 239 -37
rect 145 -71 163 -54
rect 93 -109 163 -71
rect 221 -71 239 -54
rect 273 -54 289 -37
rect 351 -37 417 -21
rect 351 -54 367 -37
rect 273 -71 291 -54
rect 221 -109 291 -71
rect 349 -71 367 -54
rect 401 -54 417 -37
rect 479 -37 545 -21
rect 479 -54 495 -37
rect 401 -71 419 -54
rect 349 -109 419 -71
rect 477 -71 495 -54
rect 529 -54 545 -37
rect 607 -37 673 -21
rect 607 -54 623 -37
rect 529 -71 547 -54
rect 477 -109 547 -71
rect 605 -71 623 -54
rect 657 -54 673 -37
rect 735 -37 801 -21
rect 735 -54 751 -37
rect 657 -71 675 -54
rect 605 -109 675 -71
rect 733 -71 751 -54
rect 785 -54 801 -37
rect 863 -37 929 -21
rect 863 -54 879 -37
rect 785 -71 803 -54
rect 733 -109 803 -71
rect 861 -71 879 -54
rect 913 -54 929 -37
rect 991 -37 1057 -21
rect 991 -54 1007 -37
rect 913 -71 931 -54
rect 861 -109 931 -71
rect 989 -71 1007 -54
rect 1041 -54 1057 -37
rect 1041 -71 1059 -54
rect 989 -109 1059 -71
rect -1059 -647 -989 -609
rect -1059 -664 -1041 -647
rect -1057 -681 -1041 -664
rect -1007 -664 -989 -647
rect -931 -647 -861 -609
rect -931 -664 -913 -647
rect -1007 -681 -991 -664
rect -1057 -697 -991 -681
rect -929 -681 -913 -664
rect -879 -664 -861 -647
rect -803 -647 -733 -609
rect -803 -664 -785 -647
rect -879 -681 -863 -664
rect -929 -697 -863 -681
rect -801 -681 -785 -664
rect -751 -664 -733 -647
rect -675 -647 -605 -609
rect -675 -664 -657 -647
rect -751 -681 -735 -664
rect -801 -697 -735 -681
rect -673 -681 -657 -664
rect -623 -664 -605 -647
rect -547 -647 -477 -609
rect -547 -664 -529 -647
rect -623 -681 -607 -664
rect -673 -697 -607 -681
rect -545 -681 -529 -664
rect -495 -664 -477 -647
rect -419 -647 -349 -609
rect -419 -664 -401 -647
rect -495 -681 -479 -664
rect -545 -697 -479 -681
rect -417 -681 -401 -664
rect -367 -664 -349 -647
rect -291 -647 -221 -609
rect -291 -664 -273 -647
rect -367 -681 -351 -664
rect -417 -697 -351 -681
rect -289 -681 -273 -664
rect -239 -664 -221 -647
rect -163 -647 -93 -609
rect -163 -664 -145 -647
rect -239 -681 -223 -664
rect -289 -697 -223 -681
rect -161 -681 -145 -664
rect -111 -664 -93 -647
rect -35 -647 35 -609
rect -35 -664 -17 -647
rect -111 -681 -95 -664
rect -161 -697 -95 -681
rect -33 -681 -17 -664
rect 17 -664 35 -647
rect 93 -647 163 -609
rect 93 -664 111 -647
rect 17 -681 33 -664
rect -33 -697 33 -681
rect 95 -681 111 -664
rect 145 -664 163 -647
rect 221 -647 291 -609
rect 221 -664 239 -647
rect 145 -681 161 -664
rect 95 -697 161 -681
rect 223 -681 239 -664
rect 273 -664 291 -647
rect 349 -647 419 -609
rect 349 -664 367 -647
rect 273 -681 289 -664
rect 223 -697 289 -681
rect 351 -681 367 -664
rect 401 -664 419 -647
rect 477 -647 547 -609
rect 477 -664 495 -647
rect 401 -681 417 -664
rect 351 -697 417 -681
rect 479 -681 495 -664
rect 529 -664 547 -647
rect 605 -647 675 -609
rect 605 -664 623 -647
rect 529 -681 545 -664
rect 479 -697 545 -681
rect 607 -681 623 -664
rect 657 -664 675 -647
rect 733 -647 803 -609
rect 733 -664 751 -647
rect 657 -681 673 -664
rect 607 -697 673 -681
rect 735 -681 751 -664
rect 785 -664 803 -647
rect 861 -647 931 -609
rect 861 -664 879 -647
rect 785 -681 801 -664
rect 735 -697 801 -681
rect 863 -681 879 -664
rect 913 -664 931 -647
rect 989 -647 1059 -609
rect 989 -664 1007 -647
rect 913 -681 929 -664
rect 863 -697 929 -681
rect 991 -681 1007 -664
rect 1041 -664 1059 -647
rect 1041 -681 1057 -664
rect 991 -697 1057 -681
<< polycont >>
rect -1041 647 -1007 681
rect -913 647 -879 681
rect -785 647 -751 681
rect -657 647 -623 681
rect -529 647 -495 681
rect -401 647 -367 681
rect -273 647 -239 681
rect -145 647 -111 681
rect -17 647 17 681
rect 111 647 145 681
rect 239 647 273 681
rect 367 647 401 681
rect 495 647 529 681
rect 623 647 657 681
rect 751 647 785 681
rect 879 647 913 681
rect 1007 647 1041 681
rect -1041 37 -1007 71
rect -913 37 -879 71
rect -785 37 -751 71
rect -657 37 -623 71
rect -529 37 -495 71
rect -401 37 -367 71
rect -273 37 -239 71
rect -145 37 -111 71
rect -17 37 17 71
rect 111 37 145 71
rect 239 37 273 71
rect 367 37 401 71
rect 495 37 529 71
rect 623 37 657 71
rect 751 37 785 71
rect 879 37 913 71
rect 1007 37 1041 71
rect -1041 -71 -1007 -37
rect -913 -71 -879 -37
rect -785 -71 -751 -37
rect -657 -71 -623 -37
rect -529 -71 -495 -37
rect -401 -71 -367 -37
rect -273 -71 -239 -37
rect -145 -71 -111 -37
rect -17 -71 17 -37
rect 111 -71 145 -37
rect 239 -71 273 -37
rect 367 -71 401 -37
rect 495 -71 529 -37
rect 623 -71 657 -37
rect 751 -71 785 -37
rect 879 -71 913 -37
rect 1007 -71 1041 -37
rect -1041 -681 -1007 -647
rect -913 -681 -879 -647
rect -785 -681 -751 -647
rect -657 -681 -623 -647
rect -529 -681 -495 -647
rect -401 -681 -367 -647
rect -273 -681 -239 -647
rect -145 -681 -111 -647
rect -17 -681 17 -647
rect 111 -681 145 -647
rect 239 -681 273 -647
rect 367 -681 401 -647
rect 495 -681 529 -647
rect 623 -681 657 -647
rect 751 -681 785 -647
rect 879 -681 913 -647
rect 1007 -681 1041 -647
<< locali >>
rect -1219 749 1219 783
rect -1219 524 -1185 749
rect -1057 647 -1043 681
rect -1005 647 -991 681
rect -929 647 -915 681
rect -877 647 -863 681
rect -801 647 -787 681
rect -749 647 -735 681
rect -673 647 -659 681
rect -621 647 -607 681
rect -545 647 -531 681
rect -493 647 -479 681
rect -417 647 -403 681
rect -365 647 -351 681
rect -289 647 -275 681
rect -237 647 -223 681
rect -161 647 -147 681
rect -109 647 -95 681
rect -33 647 -19 681
rect 19 647 33 681
rect 95 647 109 681
rect 147 647 161 681
rect 223 647 237 681
rect 275 647 289 681
rect 351 647 365 681
rect 403 647 417 681
rect 479 647 493 681
rect 531 647 545 681
rect 607 647 621 681
rect 659 647 673 681
rect 735 647 749 681
rect 787 647 801 681
rect 863 647 877 681
rect 915 647 929 681
rect 991 647 1005 681
rect 1043 647 1057 681
rect -1105 407 -1071 423
rect -1105 295 -1071 311
rect -977 407 -943 423
rect -977 295 -943 311
rect -849 407 -815 423
rect -849 295 -815 311
rect -721 407 -687 423
rect -721 295 -687 311
rect -593 407 -559 423
rect -593 295 -559 311
rect -465 407 -431 423
rect -465 295 -431 311
rect -337 407 -303 423
rect -337 295 -303 311
rect -209 407 -175 423
rect -209 295 -175 311
rect -81 407 -47 423
rect -81 295 -47 311
rect 47 407 81 423
rect 47 295 81 311
rect 175 407 209 423
rect 175 295 209 311
rect 303 407 337 423
rect 303 295 337 311
rect 431 407 465 423
rect 431 295 465 311
rect 559 407 593 423
rect 559 295 593 311
rect 687 407 721 423
rect 687 295 721 311
rect 815 407 849 423
rect 815 295 849 311
rect 943 407 977 423
rect 943 295 977 311
rect 1071 407 1105 423
rect 1071 295 1105 311
rect -1057 37 -1043 71
rect -1005 37 -991 71
rect -929 37 -915 71
rect -877 37 -863 71
rect -801 37 -787 71
rect -749 37 -735 71
rect -673 37 -659 71
rect -621 37 -607 71
rect -545 37 -531 71
rect -493 37 -479 71
rect -417 37 -403 71
rect -365 37 -351 71
rect -289 37 -275 71
rect -237 37 -223 71
rect -161 37 -147 71
rect -109 37 -95 71
rect -33 37 -19 71
rect 19 37 33 71
rect 95 37 109 71
rect 147 37 161 71
rect 223 37 237 71
rect 275 37 289 71
rect 351 37 365 71
rect 403 37 417 71
rect 479 37 493 71
rect 531 37 545 71
rect 607 37 621 71
rect 659 37 673 71
rect 735 37 749 71
rect 787 37 801 71
rect 863 37 877 71
rect 915 37 929 71
rect 991 37 1005 71
rect 1043 37 1057 71
rect -1057 -71 -1043 -37
rect -1005 -71 -991 -37
rect -929 -71 -915 -37
rect -877 -71 -863 -37
rect -801 -71 -787 -37
rect -749 -71 -735 -37
rect -673 -71 -659 -37
rect -621 -71 -607 -37
rect -545 -71 -531 -37
rect -493 -71 -479 -37
rect -417 -71 -403 -37
rect -365 -71 -351 -37
rect -289 -71 -275 -37
rect -237 -71 -223 -37
rect -161 -71 -147 -37
rect -109 -71 -95 -37
rect -33 -71 -19 -37
rect 19 -71 33 -37
rect 95 -71 109 -37
rect 147 -71 161 -37
rect 223 -71 237 -37
rect 275 -71 289 -37
rect 351 -71 365 -37
rect 403 -71 417 -37
rect 479 -71 493 -37
rect 531 -71 545 -37
rect 607 -71 621 -37
rect 659 -71 673 -37
rect 735 -71 749 -37
rect 787 -71 801 -37
rect 863 -71 877 -37
rect 915 -71 929 -37
rect 991 -71 1005 -37
rect 1043 -71 1057 -37
rect -1105 -311 -1071 -295
rect -1105 -423 -1071 -407
rect -977 -311 -943 -295
rect -977 -423 -943 -407
rect -849 -311 -815 -295
rect -849 -423 -815 -407
rect -721 -311 -687 -295
rect -721 -423 -687 -407
rect -593 -311 -559 -295
rect -593 -423 -559 -407
rect -465 -311 -431 -295
rect -465 -423 -431 -407
rect -337 -311 -303 -295
rect -337 -423 -303 -407
rect -209 -311 -175 -295
rect -209 -423 -175 -407
rect -81 -311 -47 -295
rect -81 -423 -47 -407
rect 47 -311 81 -295
rect 47 -423 81 -407
rect 175 -311 209 -295
rect 175 -423 209 -407
rect 303 -311 337 -295
rect 303 -423 337 -407
rect 431 -311 465 -295
rect 431 -423 465 -407
rect 559 -311 593 -295
rect 559 -423 593 -407
rect 687 -311 721 -295
rect 687 -423 721 -407
rect 815 -311 849 -295
rect 815 -423 849 -407
rect 943 -311 977 -295
rect 943 -423 977 -407
rect 1071 -311 1105 -295
rect 1071 -423 1105 -407
rect -1219 -749 -1185 -524
rect -1057 -681 -1043 -647
rect -1005 -681 -991 -647
rect -929 -681 -915 -647
rect -877 -681 -863 -647
rect -801 -681 -787 -647
rect -749 -681 -735 -647
rect -673 -681 -659 -647
rect -621 -681 -607 -647
rect -545 -681 -531 -647
rect -493 -681 -479 -647
rect -417 -681 -403 -647
rect -365 -681 -351 -647
rect -289 -681 -275 -647
rect -237 -681 -223 -647
rect -161 -681 -147 -647
rect -109 -681 -95 -647
rect -33 -681 -19 -647
rect 19 -681 33 -647
rect 95 -681 109 -647
rect 147 -681 161 -647
rect 223 -681 237 -647
rect 275 -681 289 -647
rect 351 -681 365 -647
rect 403 -681 417 -647
rect 479 -681 493 -647
rect 531 -681 545 -647
rect 607 -681 621 -647
rect 659 -681 673 -647
rect 735 -681 749 -647
rect 787 -681 801 -647
rect 863 -681 877 -647
rect 915 -681 929 -647
rect 991 -681 1005 -647
rect 1043 -681 1057 -647
rect 1185 -749 1219 749
rect -1219 -783 1219 -749
<< viali >>
rect -1043 647 -1041 681
rect -1041 647 -1007 681
rect -1007 647 -1005 681
rect -915 647 -913 681
rect -913 647 -879 681
rect -879 647 -877 681
rect -787 647 -785 681
rect -785 647 -751 681
rect -751 647 -749 681
rect -659 647 -657 681
rect -657 647 -623 681
rect -623 647 -621 681
rect -531 647 -529 681
rect -529 647 -495 681
rect -495 647 -493 681
rect -403 647 -401 681
rect -401 647 -367 681
rect -367 647 -365 681
rect -275 647 -273 681
rect -273 647 -239 681
rect -239 647 -237 681
rect -147 647 -145 681
rect -145 647 -111 681
rect -111 647 -109 681
rect -19 647 -17 681
rect -17 647 17 681
rect 17 647 19 681
rect 109 647 111 681
rect 111 647 145 681
rect 145 647 147 681
rect 237 647 239 681
rect 239 647 273 681
rect 273 647 275 681
rect 365 647 367 681
rect 367 647 401 681
rect 401 647 403 681
rect 493 647 495 681
rect 495 647 529 681
rect 529 647 531 681
rect 621 647 623 681
rect 623 647 657 681
rect 657 647 659 681
rect 749 647 751 681
rect 751 647 785 681
rect 785 647 787 681
rect 877 647 879 681
rect 879 647 913 681
rect 913 647 915 681
rect 1005 647 1007 681
rect 1007 647 1041 681
rect 1041 647 1043 681
rect -1219 481 -1185 524
rect -1219 -481 -1185 481
rect -1105 323 -1071 395
rect -977 323 -943 395
rect -849 323 -815 395
rect -721 323 -687 395
rect -593 323 -559 395
rect -465 323 -431 395
rect -337 323 -303 395
rect -209 323 -175 395
rect -81 323 -47 395
rect 47 323 81 395
rect 175 323 209 395
rect 303 323 337 395
rect 431 323 465 395
rect 559 323 593 395
rect 687 323 721 395
rect 815 323 849 395
rect 943 323 977 395
rect 1071 323 1105 395
rect -1043 37 -1041 71
rect -1041 37 -1007 71
rect -1007 37 -1005 71
rect -915 37 -913 71
rect -913 37 -879 71
rect -879 37 -877 71
rect -787 37 -785 71
rect -785 37 -751 71
rect -751 37 -749 71
rect -659 37 -657 71
rect -657 37 -623 71
rect -623 37 -621 71
rect -531 37 -529 71
rect -529 37 -495 71
rect -495 37 -493 71
rect -403 37 -401 71
rect -401 37 -367 71
rect -367 37 -365 71
rect -275 37 -273 71
rect -273 37 -239 71
rect -239 37 -237 71
rect -147 37 -145 71
rect -145 37 -111 71
rect -111 37 -109 71
rect -19 37 -17 71
rect -17 37 17 71
rect 17 37 19 71
rect 109 37 111 71
rect 111 37 145 71
rect 145 37 147 71
rect 237 37 239 71
rect 239 37 273 71
rect 273 37 275 71
rect 365 37 367 71
rect 367 37 401 71
rect 401 37 403 71
rect 493 37 495 71
rect 495 37 529 71
rect 529 37 531 71
rect 621 37 623 71
rect 623 37 657 71
rect 657 37 659 71
rect 749 37 751 71
rect 751 37 785 71
rect 785 37 787 71
rect 877 37 879 71
rect 879 37 913 71
rect 913 37 915 71
rect 1005 37 1007 71
rect 1007 37 1041 71
rect 1041 37 1043 71
rect -1043 -71 -1041 -37
rect -1041 -71 -1007 -37
rect -1007 -71 -1005 -37
rect -915 -71 -913 -37
rect -913 -71 -879 -37
rect -879 -71 -877 -37
rect -787 -71 -785 -37
rect -785 -71 -751 -37
rect -751 -71 -749 -37
rect -659 -71 -657 -37
rect -657 -71 -623 -37
rect -623 -71 -621 -37
rect -531 -71 -529 -37
rect -529 -71 -495 -37
rect -495 -71 -493 -37
rect -403 -71 -401 -37
rect -401 -71 -367 -37
rect -367 -71 -365 -37
rect -275 -71 -273 -37
rect -273 -71 -239 -37
rect -239 -71 -237 -37
rect -147 -71 -145 -37
rect -145 -71 -111 -37
rect -111 -71 -109 -37
rect -19 -71 -17 -37
rect -17 -71 17 -37
rect 17 -71 19 -37
rect 109 -71 111 -37
rect 111 -71 145 -37
rect 145 -71 147 -37
rect 237 -71 239 -37
rect 239 -71 273 -37
rect 273 -71 275 -37
rect 365 -71 367 -37
rect 367 -71 401 -37
rect 401 -71 403 -37
rect 493 -71 495 -37
rect 495 -71 529 -37
rect 529 -71 531 -37
rect 621 -71 623 -37
rect 623 -71 657 -37
rect 657 -71 659 -37
rect 749 -71 751 -37
rect 751 -71 785 -37
rect 785 -71 787 -37
rect 877 -71 879 -37
rect 879 -71 913 -37
rect 913 -71 915 -37
rect 1005 -71 1007 -37
rect 1007 -71 1041 -37
rect 1041 -71 1043 -37
rect -1105 -395 -1071 -323
rect -977 -395 -943 -323
rect -849 -395 -815 -323
rect -721 -395 -687 -323
rect -593 -395 -559 -323
rect -465 -395 -431 -323
rect -337 -395 -303 -323
rect -209 -395 -175 -323
rect -81 -395 -47 -323
rect 47 -395 81 -323
rect 175 -395 209 -323
rect 303 -395 337 -323
rect 431 -395 465 -323
rect 559 -395 593 -323
rect 687 -395 721 -323
rect 815 -395 849 -323
rect 943 -395 977 -323
rect 1071 -395 1105 -323
rect -1219 -524 -1185 -481
rect -1043 -681 -1041 -647
rect -1041 -681 -1007 -647
rect -1007 -681 -1005 -647
rect -915 -681 -913 -647
rect -913 -681 -879 -647
rect -879 -681 -877 -647
rect -787 -681 -785 -647
rect -785 -681 -751 -647
rect -751 -681 -749 -647
rect -659 -681 -657 -647
rect -657 -681 -623 -647
rect -623 -681 -621 -647
rect -531 -681 -529 -647
rect -529 -681 -495 -647
rect -495 -681 -493 -647
rect -403 -681 -401 -647
rect -401 -681 -367 -647
rect -367 -681 -365 -647
rect -275 -681 -273 -647
rect -273 -681 -239 -647
rect -239 -681 -237 -647
rect -147 -681 -145 -647
rect -145 -681 -111 -647
rect -111 -681 -109 -647
rect -19 -681 -17 -647
rect -17 -681 17 -647
rect 17 -681 19 -647
rect 109 -681 111 -647
rect 111 -681 145 -647
rect 145 -681 147 -647
rect 237 -681 239 -647
rect 239 -681 273 -647
rect 273 -681 275 -647
rect 365 -681 367 -647
rect 367 -681 401 -647
rect 401 -681 403 -647
rect 493 -681 495 -647
rect 495 -681 529 -647
rect 529 -681 531 -647
rect 621 -681 623 -647
rect 623 -681 657 -647
rect 657 -681 659 -647
rect 749 -681 751 -647
rect 751 -681 785 -647
rect 785 -681 787 -647
rect 877 -681 879 -647
rect 879 -681 913 -647
rect 913 -681 915 -647
rect 1005 -681 1007 -647
rect 1007 -681 1041 -647
rect 1041 -681 1043 -647
<< metal1 >>
rect -1055 681 -993 687
rect -1055 647 -1043 681
rect -1005 647 -993 681
rect -1055 641 -993 647
rect -927 681 -865 687
rect -927 647 -915 681
rect -877 647 -865 681
rect -927 641 -865 647
rect -799 681 -737 687
rect -799 647 -787 681
rect -749 647 -737 681
rect -799 641 -737 647
rect -671 681 -609 687
rect -671 647 -659 681
rect -621 647 -609 681
rect -671 641 -609 647
rect -543 681 -481 687
rect -543 647 -531 681
rect -493 647 -481 681
rect -543 641 -481 647
rect -415 681 -353 687
rect -415 647 -403 681
rect -365 647 -353 681
rect -415 641 -353 647
rect -287 681 -225 687
rect -287 647 -275 681
rect -237 647 -225 681
rect -287 641 -225 647
rect -159 681 -97 687
rect -159 647 -147 681
rect -109 647 -97 681
rect -159 641 -97 647
rect -31 681 31 687
rect -31 647 -19 681
rect 19 647 31 681
rect -31 641 31 647
rect 97 681 159 687
rect 97 647 109 681
rect 147 647 159 681
rect 97 641 159 647
rect 225 681 287 687
rect 225 647 237 681
rect 275 647 287 681
rect 225 641 287 647
rect 353 681 415 687
rect 353 647 365 681
rect 403 647 415 681
rect 353 641 415 647
rect 481 681 543 687
rect 481 647 493 681
rect 531 647 543 681
rect 481 641 543 647
rect 609 681 671 687
rect 609 647 621 681
rect 659 647 671 681
rect 609 641 671 647
rect 737 681 799 687
rect 737 647 749 681
rect 787 647 799 681
rect 737 641 799 647
rect 865 681 927 687
rect 865 647 877 681
rect 915 647 927 681
rect 865 641 927 647
rect 993 681 1055 687
rect 993 647 1005 681
rect 1043 647 1055 681
rect 993 641 1055 647
rect -1225 524 -1179 536
rect -1225 -524 -1219 524
rect -1185 -524 -1179 524
rect -1111 395 -1065 407
rect -1111 323 -1105 395
rect -1071 323 -1065 395
rect -1111 311 -1065 323
rect -983 395 -937 407
rect -983 323 -977 395
rect -943 323 -937 395
rect -983 311 -937 323
rect -855 395 -809 407
rect -855 323 -849 395
rect -815 323 -809 395
rect -855 311 -809 323
rect -727 395 -681 407
rect -727 323 -721 395
rect -687 323 -681 395
rect -727 311 -681 323
rect -599 395 -553 407
rect -599 323 -593 395
rect -559 323 -553 395
rect -599 311 -553 323
rect -471 395 -425 407
rect -471 323 -465 395
rect -431 323 -425 395
rect -471 311 -425 323
rect -343 395 -297 407
rect -343 323 -337 395
rect -303 323 -297 395
rect -343 311 -297 323
rect -215 395 -169 407
rect -215 323 -209 395
rect -175 323 -169 395
rect -215 311 -169 323
rect -87 395 -41 407
rect -87 323 -81 395
rect -47 323 -41 395
rect -87 311 -41 323
rect 41 395 87 407
rect 41 323 47 395
rect 81 323 87 395
rect 41 311 87 323
rect 169 395 215 407
rect 169 323 175 395
rect 209 323 215 395
rect 169 311 215 323
rect 297 395 343 407
rect 297 323 303 395
rect 337 323 343 395
rect 297 311 343 323
rect 425 395 471 407
rect 425 323 431 395
rect 465 323 471 395
rect 425 311 471 323
rect 553 395 599 407
rect 553 323 559 395
rect 593 323 599 395
rect 553 311 599 323
rect 681 395 727 407
rect 681 323 687 395
rect 721 323 727 395
rect 681 311 727 323
rect 809 395 855 407
rect 809 323 815 395
rect 849 323 855 395
rect 809 311 855 323
rect 937 395 983 407
rect 937 323 943 395
rect 977 323 983 395
rect 937 311 983 323
rect 1065 395 1111 407
rect 1065 323 1071 395
rect 1105 323 1111 395
rect 1065 311 1111 323
rect -1055 71 -993 77
rect -1055 37 -1043 71
rect -1005 37 -993 71
rect -1055 31 -993 37
rect -927 71 -865 77
rect -927 37 -915 71
rect -877 37 -865 71
rect -927 31 -865 37
rect -799 71 -737 77
rect -799 37 -787 71
rect -749 37 -737 71
rect -799 31 -737 37
rect -671 71 -609 77
rect -671 37 -659 71
rect -621 37 -609 71
rect -671 31 -609 37
rect -543 71 -481 77
rect -543 37 -531 71
rect -493 37 -481 71
rect -543 31 -481 37
rect -415 71 -353 77
rect -415 37 -403 71
rect -365 37 -353 71
rect -415 31 -353 37
rect -287 71 -225 77
rect -287 37 -275 71
rect -237 37 -225 71
rect -287 31 -225 37
rect -159 71 -97 77
rect -159 37 -147 71
rect -109 37 -97 71
rect -159 31 -97 37
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect 97 71 159 77
rect 97 37 109 71
rect 147 37 159 71
rect 97 31 159 37
rect 225 71 287 77
rect 225 37 237 71
rect 275 37 287 71
rect 225 31 287 37
rect 353 71 415 77
rect 353 37 365 71
rect 403 37 415 71
rect 353 31 415 37
rect 481 71 543 77
rect 481 37 493 71
rect 531 37 543 71
rect 481 31 543 37
rect 609 71 671 77
rect 609 37 621 71
rect 659 37 671 71
rect 609 31 671 37
rect 737 71 799 77
rect 737 37 749 71
rect 787 37 799 71
rect 737 31 799 37
rect 865 71 927 77
rect 865 37 877 71
rect 915 37 927 71
rect 865 31 927 37
rect 993 71 1055 77
rect 993 37 1005 71
rect 1043 37 1055 71
rect 993 31 1055 37
rect -1055 -37 -993 -31
rect -1055 -71 -1043 -37
rect -1005 -71 -993 -37
rect -1055 -77 -993 -71
rect -927 -37 -865 -31
rect -927 -71 -915 -37
rect -877 -71 -865 -37
rect -927 -77 -865 -71
rect -799 -37 -737 -31
rect -799 -71 -787 -37
rect -749 -71 -737 -37
rect -799 -77 -737 -71
rect -671 -37 -609 -31
rect -671 -71 -659 -37
rect -621 -71 -609 -37
rect -671 -77 -609 -71
rect -543 -37 -481 -31
rect -543 -71 -531 -37
rect -493 -71 -481 -37
rect -543 -77 -481 -71
rect -415 -37 -353 -31
rect -415 -71 -403 -37
rect -365 -71 -353 -37
rect -415 -77 -353 -71
rect -287 -37 -225 -31
rect -287 -71 -275 -37
rect -237 -71 -225 -37
rect -287 -77 -225 -71
rect -159 -37 -97 -31
rect -159 -71 -147 -37
rect -109 -71 -97 -37
rect -159 -77 -97 -71
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect 97 -37 159 -31
rect 97 -71 109 -37
rect 147 -71 159 -37
rect 97 -77 159 -71
rect 225 -37 287 -31
rect 225 -71 237 -37
rect 275 -71 287 -37
rect 225 -77 287 -71
rect 353 -37 415 -31
rect 353 -71 365 -37
rect 403 -71 415 -37
rect 353 -77 415 -71
rect 481 -37 543 -31
rect 481 -71 493 -37
rect 531 -71 543 -37
rect 481 -77 543 -71
rect 609 -37 671 -31
rect 609 -71 621 -37
rect 659 -71 671 -37
rect 609 -77 671 -71
rect 737 -37 799 -31
rect 737 -71 749 -37
rect 787 -71 799 -37
rect 737 -77 799 -71
rect 865 -37 927 -31
rect 865 -71 877 -37
rect 915 -71 927 -37
rect 865 -77 927 -71
rect 993 -37 1055 -31
rect 993 -71 1005 -37
rect 1043 -71 1055 -37
rect 993 -77 1055 -71
rect -1111 -323 -1065 -311
rect -1111 -395 -1105 -323
rect -1071 -395 -1065 -323
rect -1111 -407 -1065 -395
rect -983 -323 -937 -311
rect -983 -395 -977 -323
rect -943 -395 -937 -323
rect -983 -407 -937 -395
rect -855 -323 -809 -311
rect -855 -395 -849 -323
rect -815 -395 -809 -323
rect -855 -407 -809 -395
rect -727 -323 -681 -311
rect -727 -395 -721 -323
rect -687 -395 -681 -323
rect -727 -407 -681 -395
rect -599 -323 -553 -311
rect -599 -395 -593 -323
rect -559 -395 -553 -323
rect -599 -407 -553 -395
rect -471 -323 -425 -311
rect -471 -395 -465 -323
rect -431 -395 -425 -323
rect -471 -407 -425 -395
rect -343 -323 -297 -311
rect -343 -395 -337 -323
rect -303 -395 -297 -323
rect -343 -407 -297 -395
rect -215 -323 -169 -311
rect -215 -395 -209 -323
rect -175 -395 -169 -323
rect -215 -407 -169 -395
rect -87 -323 -41 -311
rect -87 -395 -81 -323
rect -47 -395 -41 -323
rect -87 -407 -41 -395
rect 41 -323 87 -311
rect 41 -395 47 -323
rect 81 -395 87 -323
rect 41 -407 87 -395
rect 169 -323 215 -311
rect 169 -395 175 -323
rect 209 -395 215 -323
rect 169 -407 215 -395
rect 297 -323 343 -311
rect 297 -395 303 -323
rect 337 -395 343 -323
rect 297 -407 343 -395
rect 425 -323 471 -311
rect 425 -395 431 -323
rect 465 -395 471 -323
rect 425 -407 471 -395
rect 553 -323 599 -311
rect 553 -395 559 -323
rect 593 -395 599 -323
rect 553 -407 599 -395
rect 681 -323 727 -311
rect 681 -395 687 -323
rect 721 -395 727 -323
rect 681 -407 727 -395
rect 809 -323 855 -311
rect 809 -395 815 -323
rect 849 -395 855 -323
rect 809 -407 855 -395
rect 937 -323 983 -311
rect 937 -395 943 -323
rect 977 -395 983 -323
rect 937 -407 983 -395
rect 1065 -323 1111 -311
rect 1065 -395 1071 -323
rect 1105 -395 1111 -323
rect 1065 -407 1111 -395
rect -1225 -536 -1179 -524
rect -1055 -647 -993 -641
rect -1055 -681 -1043 -647
rect -1005 -681 -993 -647
rect -1055 -687 -993 -681
rect -927 -647 -865 -641
rect -927 -681 -915 -647
rect -877 -681 -865 -647
rect -927 -687 -865 -681
rect -799 -647 -737 -641
rect -799 -681 -787 -647
rect -749 -681 -737 -647
rect -799 -687 -737 -681
rect -671 -647 -609 -641
rect -671 -681 -659 -647
rect -621 -681 -609 -647
rect -671 -687 -609 -681
rect -543 -647 -481 -641
rect -543 -681 -531 -647
rect -493 -681 -481 -647
rect -543 -687 -481 -681
rect -415 -647 -353 -641
rect -415 -681 -403 -647
rect -365 -681 -353 -647
rect -415 -687 -353 -681
rect -287 -647 -225 -641
rect -287 -681 -275 -647
rect -237 -681 -225 -647
rect -287 -687 -225 -681
rect -159 -647 -97 -641
rect -159 -681 -147 -647
rect -109 -681 -97 -647
rect -159 -687 -97 -681
rect -31 -647 31 -641
rect -31 -681 -19 -647
rect 19 -681 31 -647
rect -31 -687 31 -681
rect 97 -647 159 -641
rect 97 -681 109 -647
rect 147 -681 159 -647
rect 97 -687 159 -681
rect 225 -647 287 -641
rect 225 -681 237 -647
rect 275 -681 287 -647
rect 225 -687 287 -681
rect 353 -647 415 -641
rect 353 -681 365 -647
rect 403 -681 415 -647
rect 353 -687 415 -681
rect 481 -647 543 -641
rect 481 -681 493 -647
rect 531 -681 543 -647
rect 481 -687 543 -681
rect 609 -647 671 -641
rect 609 -681 621 -647
rect 659 -681 671 -647
rect 609 -687 671 -681
rect 737 -647 799 -641
rect 737 -681 749 -647
rect 787 -681 799 -647
rect 737 -687 799 -681
rect 865 -647 927 -641
rect 865 -681 877 -647
rect 915 -681 927 -647
rect 865 -687 927 -681
rect 993 -647 1055 -641
rect 993 -681 1005 -647
rect 1043 -681 1055 -647
rect 993 -687 1055 -681
<< properties >>
string FIXED_BBOX -1202 -766 1202 766
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.5 l 0.35 m 2 nf 17 diffcov 20 polycov 70 guard 1 glc 1 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 15 viadrn 15 viagate 100 viagb 0 viagr 0 viagl 70 viagt 0
<< end >>
