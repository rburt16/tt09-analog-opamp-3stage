magic
tech sky130A
magscale 1 2
timestamp 1730569394
<< nwell >>
rect -554 -1219 554 1219
<< pmos >>
rect -358 -1000 -158 1000
rect -100 -1000 100 1000
rect 158 -1000 358 1000
<< pdiff >>
rect -416 692 -358 1000
rect -416 -692 -404 692
rect -370 -692 -358 692
rect -416 -1000 -358 -692
rect -158 692 -100 1000
rect -158 -692 -146 692
rect -112 -692 -100 692
rect -158 -1000 -100 -692
rect 100 692 158 1000
rect 100 -692 112 692
rect 146 -692 158 692
rect 100 -1000 158 -692
rect 358 692 416 1000
rect 358 -692 370 692
rect 404 -692 416 692
rect 358 -1000 416 -692
<< pdiffc >>
rect -404 -692 -370 692
rect -146 -692 -112 692
rect 112 -692 146 692
rect 370 -692 404 692
<< nsubdiff >>
rect -518 1149 -295 1183
rect 295 1149 518 1183
rect -518 761 -484 1149
rect -518 -1149 -484 -761
rect 484 761 518 1149
rect 484 -1149 518 -761
rect -518 -1183 -295 -1149
rect 295 -1183 518 -1149
<< nsubdiffcont >>
rect -295 1149 295 1183
rect -518 -761 -484 761
rect 484 -761 518 761
rect -295 -1183 295 -1149
<< poly >>
rect -333 1081 -183 1097
rect -333 1064 -317 1081
rect -358 1047 -317 1064
rect -199 1064 -183 1081
rect -75 1081 75 1097
rect -75 1064 -59 1081
rect -199 1047 -158 1064
rect -358 1000 -158 1047
rect -100 1047 -59 1064
rect 59 1064 75 1081
rect 183 1081 333 1097
rect 183 1064 199 1081
rect 59 1047 100 1064
rect -100 1000 100 1047
rect 158 1047 199 1064
rect 317 1064 333 1081
rect 317 1047 358 1064
rect 158 1000 358 1047
rect -358 -1047 -158 -1000
rect -358 -1064 -317 -1047
rect -333 -1081 -317 -1064
rect -199 -1064 -158 -1047
rect -100 -1047 100 -1000
rect -100 -1064 -59 -1047
rect -199 -1081 -183 -1064
rect -333 -1097 -183 -1081
rect -75 -1081 -59 -1064
rect 59 -1064 100 -1047
rect 158 -1047 358 -1000
rect 158 -1064 199 -1047
rect 59 -1081 75 -1064
rect -75 -1097 75 -1081
rect 183 -1081 199 -1064
rect 317 -1064 358 -1047
rect 317 -1081 333 -1064
rect 183 -1097 333 -1081
<< polycont >>
rect -317 1047 -199 1081
rect -59 1047 59 1081
rect 199 1047 317 1081
rect -317 -1081 -199 -1047
rect -59 -1081 59 -1047
rect 199 -1081 317 -1047
<< locali >>
rect -518 1149 -339 1183
rect 339 1149 518 1183
rect -518 804 -484 1149
rect 484 804 518 1149
rect -404 692 -370 708
rect -404 -708 -370 -692
rect -146 692 -112 708
rect -146 -708 -112 -692
rect 112 692 146 708
rect 112 -708 146 -692
rect 370 692 404 708
rect 370 -708 404 -692
rect -518 -1149 -484 -804
rect 484 -1149 518 -804
rect -518 -1183 -339 -1149
rect 339 -1183 518 -1149
<< viali >>
rect -339 1149 -295 1183
rect -295 1149 295 1183
rect 295 1149 339 1183
rect -342 1047 -317 1081
rect -317 1047 -199 1081
rect -199 1047 -174 1081
rect -84 1047 -59 1081
rect -59 1047 59 1081
rect 59 1047 84 1081
rect 174 1047 199 1081
rect 199 1047 317 1081
rect 317 1047 342 1081
rect -518 761 -484 804
rect -518 -761 -484 761
rect 484 761 518 804
rect -404 -692 -370 692
rect -146 -692 -112 692
rect 112 -692 146 692
rect 370 -692 404 692
rect -518 -804 -484 -761
rect 484 -761 518 761
rect 484 -804 518 -761
rect -342 -1081 -317 -1047
rect -317 -1081 -199 -1047
rect -199 -1081 -174 -1047
rect -84 -1081 -59 -1047
rect -59 -1081 59 -1047
rect 59 -1081 84 -1047
rect 174 -1081 199 -1047
rect 199 -1081 317 -1047
rect 317 -1081 342 -1047
rect -339 -1183 -295 -1149
rect -295 -1183 295 -1149
rect 295 -1183 339 -1149
<< metal1 >>
rect -351 1183 351 1189
rect -351 1149 -339 1183
rect 339 1149 351 1183
rect -351 1143 351 1149
rect -354 1081 -162 1087
rect -354 1047 -342 1081
rect -174 1047 -162 1081
rect -354 1041 -162 1047
rect -96 1081 96 1087
rect -96 1047 -84 1081
rect 84 1047 96 1081
rect -96 1041 96 1047
rect 162 1081 354 1087
rect 162 1047 174 1081
rect 342 1047 354 1081
rect 162 1041 354 1047
rect -524 804 -478 816
rect -524 -804 -518 804
rect -484 -804 -478 804
rect 478 804 524 816
rect -410 692 -364 704
rect -410 -692 -404 692
rect -370 -692 -364 692
rect -410 -704 -364 -692
rect -152 692 -106 704
rect -152 -692 -146 692
rect -112 -692 -106 692
rect -152 -704 -106 -692
rect 106 692 152 704
rect 106 -692 112 692
rect 146 -692 152 692
rect 106 -704 152 -692
rect 364 692 410 704
rect 364 -692 370 692
rect 404 -692 410 692
rect 364 -704 410 -692
rect -524 -816 -478 -804
rect 478 -804 484 804
rect 518 -804 524 804
rect 478 -816 524 -804
rect -354 -1047 -162 -1041
rect -354 -1081 -342 -1047
rect -174 -1081 -162 -1047
rect -354 -1087 -162 -1081
rect -96 -1047 96 -1041
rect -96 -1081 -84 -1047
rect 84 -1081 96 -1047
rect -96 -1087 96 -1081
rect 162 -1047 354 -1041
rect 162 -1081 174 -1047
rect 342 -1081 354 -1047
rect 162 -1087 354 -1081
rect -351 -1149 351 -1143
rect -351 -1183 -339 -1149
rect 339 -1183 351 -1149
rect -351 -1189 351 -1183
<< properties >>
string FIXED_BBOX -501 -1166 501 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 1 nf 3 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
