VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rburt16_opamp_3stage
  CLASS BLOCK ;
  FOREIGN tt_um_rburt16_opamp_3stage ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 47.849998 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 896.000000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 896.000000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.375000 ;
    ANTENNADIFFAREA 261.713989 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.750 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.750 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 12.000 177.650 17.540 189.840 ;
        RECT 18.850 177.650 21.160 189.840 ;
        RECT 12.000 130.650 17.540 176.380 ;
        RECT 18.850 130.650 21.160 176.380 ;
        RECT 22.450 130.800 27.990 176.530 ;
        RECT 29.300 130.800 31.610 176.530 ;
        RECT 32.900 159.900 38.440 183.270 ;
        RECT 39.750 159.900 42.060 183.270 ;
        RECT 43.350 159.900 48.890 183.270 ;
        RECT 50.200 159.900 52.510 183.270 ;
        RECT 60.250 177.550 62.560 189.740 ;
        RECT 63.850 177.550 66.160 189.740 ;
        RECT 67.450 177.550 69.760 189.740 ;
        RECT 74.450 166.350 83.160 189.720 ;
      LAYER pwell ;
        RECT 60.200 161.150 62.510 165.750 ;
        RECT 63.800 161.150 66.110 165.750 ;
        RECT 67.450 161.200 69.760 165.800 ;
        RECT 34.850 139.450 40.810 158.640 ;
      LAYER nwell ;
        RECT 12.000 117.150 17.540 129.340 ;
        RECT 18.850 117.150 21.160 129.340 ;
        RECT 22.450 117.300 27.990 129.490 ;
        RECT 29.300 117.300 31.610 129.490 ;
      LAYER pwell ;
        RECT 32.050 128.600 34.360 133.200 ;
        RECT 34.850 128.600 40.810 138.700 ;
        RECT 32.050 117.750 34.360 122.350 ;
        RECT 34.855 117.755 40.815 127.855 ;
        RECT 45.450 117.000 51.410 158.910 ;
        RECT 72.550 157.600 85.100 165.790 ;
        RECT 75.000 146.250 77.960 150.040 ;
        RECT 79.250 146.250 82.210 150.040 ;
      LAYER nwell ;
        RECT 22.950 115.840 25.910 115.845 ;
        RECT 12.120 106.000 17.510 115.840 ;
      LAYER pwell ;
        RECT 17.520 106.000 20.480 115.790 ;
      LAYER nwell ;
        RECT 20.520 106.005 25.910 115.840 ;
      LAYER pwell ;
        RECT 25.930 106.015 28.890 115.805 ;
      LAYER nwell ;
        RECT 28.920 111.260 39.075 115.840 ;
      LAYER pwell ;
        RECT 39.120 111.300 49.080 113.510 ;
      LAYER nwell ;
        RECT 28.920 109.000 48.580 111.260 ;
        RECT 20.520 106.000 23.480 106.005 ;
        RECT 28.920 106.000 39.075 109.000 ;
      LAYER pwell ;
        RECT 39.120 106.000 48.910 108.960 ;
        RECT 12.100 105.590 34.500 105.690 ;
        RECT 12.100 102.800 49.080 105.590 ;
        RECT 12.100 95.900 43.980 102.800 ;
        RECT 53.100 93.200 59.060 135.110 ;
      LAYER nwell ;
        RECT 74.300 133.150 77.950 145.340 ;
        RECT 79.250 133.150 82.900 145.340 ;
      LAYER pwell ;
        RECT 59.700 109.850 77.950 131.950 ;
        RECT 79.250 109.850 97.500 131.950 ;
      LAYER nwell ;
        RECT 98.250 118.100 100.560 130.290 ;
        RECT 101.850 118.100 104.160 130.290 ;
        RECT 105.450 118.100 107.760 130.290 ;
        RECT 109.050 118.100 111.360 122.790 ;
      LAYER pwell ;
        RECT 46.700 85.450 52.660 90.550 ;
        RECT 53.100 85.450 59.060 90.550 ;
        RECT 59.700 86.450 77.950 108.550 ;
        RECT 79.250 86.450 97.500 108.550 ;
        RECT 98.250 95.500 116.500 117.600 ;
      LAYER nwell ;
        RECT 44.600 62.950 77.950 85.140 ;
        RECT 79.250 62.950 112.600 85.140 ;
        RECT 44.600 39.450 77.950 61.640 ;
        RECT 79.250 39.450 112.600 61.640 ;
      LAYER li1 ;
        RECT 12.180 189.490 17.360 189.660 ;
        RECT 12.180 178.000 12.350 189.490 ;
        RECT 13.060 188.980 13.900 189.150 ;
        RECT 14.350 188.980 15.190 189.150 ;
        RECT 15.640 188.980 16.480 189.150 ;
        RECT 12.750 180.205 12.920 187.285 ;
        RECT 14.040 180.205 14.210 187.285 ;
        RECT 15.330 180.205 15.500 187.285 ;
        RECT 16.620 180.205 16.790 187.285 ;
        RECT 13.060 178.340 13.900 178.510 ;
        RECT 14.350 178.340 15.190 178.510 ;
        RECT 15.640 178.340 16.480 178.510 ;
        RECT 17.190 178.000 17.360 189.490 ;
        RECT 12.180 177.830 17.360 178.000 ;
        RECT 19.030 189.490 20.980 189.660 ;
        RECT 19.030 178.000 19.200 189.490 ;
        RECT 19.840 188.980 20.170 189.150 ;
        RECT 19.600 180.205 19.770 187.285 ;
        RECT 20.240 180.205 20.410 187.285 ;
        RECT 19.840 178.340 20.170 178.510 ;
        RECT 20.810 178.000 20.980 189.490 ;
        RECT 60.430 189.390 62.380 189.560 ;
        RECT 19.030 177.830 20.980 178.000 ;
        RECT 33.080 182.920 38.260 183.090 ;
        RECT 12.180 176.030 17.360 176.200 ;
        RECT 12.180 131.000 12.350 176.030 ;
        RECT 13.060 175.520 13.900 175.690 ;
        RECT 14.350 175.520 15.190 175.690 ;
        RECT 15.640 175.520 16.480 175.690 ;
        RECT 12.750 166.745 12.920 173.825 ;
        RECT 14.040 166.745 14.210 173.825 ;
        RECT 15.330 166.745 15.500 173.825 ;
        RECT 16.620 166.745 16.790 173.825 ;
        RECT 13.060 164.880 13.900 165.050 ;
        RECT 14.350 164.880 15.190 165.050 ;
        RECT 15.640 164.880 16.480 165.050 ;
        RECT 13.060 164.340 13.900 164.510 ;
        RECT 14.350 164.340 15.190 164.510 ;
        RECT 15.640 164.340 16.480 164.510 ;
        RECT 12.750 155.565 12.920 162.645 ;
        RECT 14.040 155.565 14.210 162.645 ;
        RECT 15.330 155.565 15.500 162.645 ;
        RECT 16.620 155.565 16.790 162.645 ;
        RECT 13.060 153.700 13.900 153.870 ;
        RECT 14.350 153.700 15.190 153.870 ;
        RECT 15.640 153.700 16.480 153.870 ;
        RECT 13.060 153.160 13.900 153.330 ;
        RECT 14.350 153.160 15.190 153.330 ;
        RECT 15.640 153.160 16.480 153.330 ;
        RECT 12.750 144.385 12.920 151.465 ;
        RECT 14.040 144.385 14.210 151.465 ;
        RECT 15.330 144.385 15.500 151.465 ;
        RECT 16.620 144.385 16.790 151.465 ;
        RECT 13.060 142.520 13.900 142.690 ;
        RECT 14.350 142.520 15.190 142.690 ;
        RECT 15.640 142.520 16.480 142.690 ;
        RECT 13.060 141.980 13.900 142.150 ;
        RECT 14.350 141.980 15.190 142.150 ;
        RECT 15.640 141.980 16.480 142.150 ;
        RECT 12.750 133.205 12.920 140.285 ;
        RECT 14.040 133.205 14.210 140.285 ;
        RECT 15.330 133.205 15.500 140.285 ;
        RECT 16.620 133.205 16.790 140.285 ;
        RECT 13.060 131.340 13.900 131.510 ;
        RECT 14.350 131.340 15.190 131.510 ;
        RECT 15.640 131.340 16.480 131.510 ;
        RECT 17.190 131.000 17.360 176.030 ;
        RECT 12.180 130.830 17.360 131.000 ;
        RECT 19.030 176.030 20.980 176.200 ;
        RECT 19.030 131.000 19.200 176.030 ;
        RECT 19.840 175.520 20.170 175.690 ;
        RECT 19.600 166.745 19.770 173.825 ;
        RECT 20.240 166.745 20.410 173.825 ;
        RECT 19.840 164.880 20.170 165.050 ;
        RECT 19.840 164.340 20.170 164.510 ;
        RECT 19.600 155.565 19.770 162.645 ;
        RECT 20.240 155.565 20.410 162.645 ;
        RECT 19.840 153.700 20.170 153.870 ;
        RECT 19.840 153.160 20.170 153.330 ;
        RECT 19.600 144.385 19.770 151.465 ;
        RECT 20.240 144.385 20.410 151.465 ;
        RECT 19.840 142.520 20.170 142.690 ;
        RECT 19.840 141.980 20.170 142.150 ;
        RECT 19.600 133.205 19.770 140.285 ;
        RECT 20.240 133.205 20.410 140.285 ;
        RECT 19.840 131.340 20.170 131.510 ;
        RECT 20.810 131.000 20.980 176.030 ;
        RECT 19.030 130.830 20.980 131.000 ;
        RECT 22.630 176.180 27.810 176.350 ;
        RECT 22.630 131.150 22.800 176.180 ;
        RECT 23.510 175.670 24.350 175.840 ;
        RECT 24.800 175.670 25.640 175.840 ;
        RECT 26.090 175.670 26.930 175.840 ;
        RECT 23.200 166.895 23.370 173.975 ;
        RECT 24.490 166.895 24.660 173.975 ;
        RECT 25.780 166.895 25.950 173.975 ;
        RECT 27.070 166.895 27.240 173.975 ;
        RECT 23.510 165.030 24.350 165.200 ;
        RECT 24.800 165.030 25.640 165.200 ;
        RECT 26.090 165.030 26.930 165.200 ;
        RECT 23.510 164.490 24.350 164.660 ;
        RECT 24.800 164.490 25.640 164.660 ;
        RECT 26.090 164.490 26.930 164.660 ;
        RECT 23.200 155.715 23.370 162.795 ;
        RECT 24.490 155.715 24.660 162.795 ;
        RECT 25.780 155.715 25.950 162.795 ;
        RECT 27.070 155.715 27.240 162.795 ;
        RECT 23.510 153.850 24.350 154.020 ;
        RECT 24.800 153.850 25.640 154.020 ;
        RECT 26.090 153.850 26.930 154.020 ;
        RECT 23.510 153.310 24.350 153.480 ;
        RECT 24.800 153.310 25.640 153.480 ;
        RECT 26.090 153.310 26.930 153.480 ;
        RECT 23.200 144.535 23.370 151.615 ;
        RECT 24.490 144.535 24.660 151.615 ;
        RECT 25.780 144.535 25.950 151.615 ;
        RECT 27.070 144.535 27.240 151.615 ;
        RECT 23.510 142.670 24.350 142.840 ;
        RECT 24.800 142.670 25.640 142.840 ;
        RECT 26.090 142.670 26.930 142.840 ;
        RECT 23.510 142.130 24.350 142.300 ;
        RECT 24.800 142.130 25.640 142.300 ;
        RECT 26.090 142.130 26.930 142.300 ;
        RECT 23.200 133.355 23.370 140.435 ;
        RECT 24.490 133.355 24.660 140.435 ;
        RECT 25.780 133.355 25.950 140.435 ;
        RECT 27.070 133.355 27.240 140.435 ;
        RECT 23.510 131.490 24.350 131.660 ;
        RECT 24.800 131.490 25.640 131.660 ;
        RECT 26.090 131.490 26.930 131.660 ;
        RECT 27.640 131.150 27.810 176.180 ;
        RECT 22.630 130.980 27.810 131.150 ;
        RECT 29.480 176.180 31.430 176.350 ;
        RECT 29.480 131.150 29.650 176.180 ;
        RECT 30.290 175.670 30.620 175.840 ;
        RECT 30.050 166.895 30.220 173.975 ;
        RECT 30.690 166.895 30.860 173.975 ;
        RECT 30.290 165.030 30.620 165.200 ;
        RECT 30.290 164.490 30.620 164.660 ;
        RECT 30.050 155.715 30.220 162.795 ;
        RECT 30.690 155.715 30.860 162.795 ;
        RECT 30.290 153.850 30.620 154.020 ;
        RECT 30.290 153.310 30.620 153.480 ;
        RECT 30.050 144.535 30.220 151.615 ;
        RECT 30.690 144.535 30.860 151.615 ;
        RECT 30.290 142.670 30.620 142.840 ;
        RECT 30.290 142.130 30.620 142.300 ;
        RECT 30.050 133.355 30.220 140.435 ;
        RECT 30.690 133.355 30.860 140.435 ;
        RECT 30.290 131.490 30.620 131.660 ;
        RECT 31.260 131.150 31.430 176.180 ;
        RECT 33.080 160.250 33.250 182.920 ;
        RECT 33.960 182.410 34.800 182.580 ;
        RECT 35.250 182.410 36.090 182.580 ;
        RECT 36.540 182.410 37.380 182.580 ;
        RECT 33.650 173.635 33.820 180.715 ;
        RECT 34.940 173.635 35.110 180.715 ;
        RECT 36.230 173.635 36.400 180.715 ;
        RECT 37.520 173.635 37.690 180.715 ;
        RECT 33.960 171.770 34.800 171.940 ;
        RECT 35.250 171.770 36.090 171.940 ;
        RECT 36.540 171.770 37.380 171.940 ;
        RECT 33.960 171.230 34.800 171.400 ;
        RECT 35.250 171.230 36.090 171.400 ;
        RECT 36.540 171.230 37.380 171.400 ;
        RECT 33.650 162.455 33.820 169.535 ;
        RECT 34.940 162.455 35.110 169.535 ;
        RECT 36.230 162.455 36.400 169.535 ;
        RECT 37.520 162.455 37.690 169.535 ;
        RECT 33.960 160.590 34.800 160.760 ;
        RECT 35.250 160.590 36.090 160.760 ;
        RECT 36.540 160.590 37.380 160.760 ;
        RECT 38.090 160.250 38.260 182.920 ;
        RECT 33.080 160.080 38.260 160.250 ;
        RECT 39.930 182.920 41.880 183.090 ;
        RECT 39.930 160.250 40.100 182.920 ;
        RECT 40.740 182.410 41.070 182.580 ;
        RECT 40.500 173.635 40.670 180.715 ;
        RECT 41.140 173.635 41.310 180.715 ;
        RECT 40.740 171.770 41.070 171.940 ;
        RECT 40.740 171.230 41.070 171.400 ;
        RECT 40.500 162.455 40.670 169.535 ;
        RECT 41.140 162.455 41.310 169.535 ;
        RECT 40.740 160.590 41.070 160.760 ;
        RECT 41.710 160.250 41.880 182.920 ;
        RECT 39.930 160.080 41.880 160.250 ;
        RECT 43.530 182.920 48.710 183.090 ;
        RECT 43.530 160.250 43.700 182.920 ;
        RECT 44.410 182.410 45.250 182.580 ;
        RECT 45.700 182.410 46.540 182.580 ;
        RECT 46.990 182.410 47.830 182.580 ;
        RECT 44.100 173.635 44.270 180.715 ;
        RECT 45.390 173.635 45.560 180.715 ;
        RECT 46.680 173.635 46.850 180.715 ;
        RECT 47.970 173.635 48.140 180.715 ;
        RECT 44.410 171.770 45.250 171.940 ;
        RECT 45.700 171.770 46.540 171.940 ;
        RECT 46.990 171.770 47.830 171.940 ;
        RECT 44.410 171.230 45.250 171.400 ;
        RECT 45.700 171.230 46.540 171.400 ;
        RECT 46.990 171.230 47.830 171.400 ;
        RECT 44.100 162.455 44.270 169.535 ;
        RECT 45.390 162.455 45.560 169.535 ;
        RECT 46.680 162.455 46.850 169.535 ;
        RECT 47.970 162.455 48.140 169.535 ;
        RECT 44.410 160.590 45.250 160.760 ;
        RECT 45.700 160.590 46.540 160.760 ;
        RECT 46.990 160.590 47.830 160.760 ;
        RECT 48.540 160.250 48.710 182.920 ;
        RECT 43.530 160.080 48.710 160.250 ;
        RECT 50.380 182.920 52.330 183.090 ;
        RECT 50.380 160.250 50.550 182.920 ;
        RECT 51.190 182.410 51.520 182.580 ;
        RECT 50.950 173.635 51.120 180.715 ;
        RECT 51.590 173.635 51.760 180.715 ;
        RECT 51.190 171.770 51.520 171.940 ;
        RECT 51.190 171.230 51.520 171.400 ;
        RECT 50.950 162.455 51.120 169.535 ;
        RECT 51.590 162.455 51.760 169.535 ;
        RECT 51.190 160.590 51.520 160.760 ;
        RECT 52.160 160.250 52.330 182.920 ;
        RECT 60.430 177.900 60.600 189.390 ;
        RECT 61.240 188.880 61.570 189.050 ;
        RECT 61.000 180.105 61.170 187.185 ;
        RECT 61.640 180.105 61.810 187.185 ;
        RECT 61.240 178.240 61.570 178.410 ;
        RECT 62.210 177.900 62.380 189.390 ;
        RECT 60.430 177.730 62.380 177.900 ;
        RECT 64.030 189.390 65.980 189.560 ;
        RECT 64.030 177.900 64.200 189.390 ;
        RECT 64.840 188.880 65.170 189.050 ;
        RECT 64.600 180.105 64.770 187.185 ;
        RECT 65.240 180.105 65.410 187.185 ;
        RECT 64.840 178.240 65.170 178.410 ;
        RECT 65.810 177.900 65.980 189.390 ;
        RECT 64.030 177.730 65.980 177.900 ;
        RECT 67.630 189.390 69.580 189.560 ;
        RECT 67.630 177.900 67.800 189.390 ;
        RECT 68.440 188.880 68.770 189.050 ;
        RECT 68.200 180.105 68.370 187.185 ;
        RECT 68.840 180.105 69.010 187.185 ;
        RECT 68.440 178.240 68.770 178.410 ;
        RECT 69.410 177.900 69.580 189.390 ;
        RECT 67.630 177.730 69.580 177.900 ;
        RECT 74.630 189.370 82.980 189.540 ;
        RECT 74.630 166.700 74.800 189.370 ;
        RECT 75.440 188.860 75.770 189.030 ;
        RECT 76.080 188.860 76.410 189.030 ;
        RECT 76.720 188.860 77.050 189.030 ;
        RECT 77.360 188.860 77.690 189.030 ;
        RECT 78.000 188.860 78.330 189.030 ;
        RECT 78.640 188.860 78.970 189.030 ;
        RECT 79.280 188.860 79.610 189.030 ;
        RECT 79.920 188.860 80.250 189.030 ;
        RECT 80.560 188.860 80.890 189.030 ;
        RECT 81.200 188.860 81.530 189.030 ;
        RECT 81.840 188.860 82.170 189.030 ;
        RECT 75.200 180.085 75.370 187.165 ;
        RECT 75.840 180.085 76.010 187.165 ;
        RECT 76.480 180.085 76.650 187.165 ;
        RECT 77.120 180.085 77.290 187.165 ;
        RECT 77.760 180.085 77.930 187.165 ;
        RECT 78.400 180.085 78.570 187.165 ;
        RECT 79.040 180.085 79.210 187.165 ;
        RECT 79.680 180.085 79.850 187.165 ;
        RECT 80.320 180.085 80.490 187.165 ;
        RECT 80.960 180.085 81.130 187.165 ;
        RECT 81.600 180.085 81.770 187.165 ;
        RECT 82.240 180.085 82.410 187.165 ;
        RECT 75.440 178.220 75.770 178.390 ;
        RECT 76.080 178.220 76.410 178.390 ;
        RECT 76.720 178.220 77.050 178.390 ;
        RECT 77.360 178.220 77.690 178.390 ;
        RECT 78.000 178.220 78.330 178.390 ;
        RECT 78.640 178.220 78.970 178.390 ;
        RECT 79.280 178.220 79.610 178.390 ;
        RECT 79.920 178.220 80.250 178.390 ;
        RECT 80.560 178.220 80.890 178.390 ;
        RECT 81.200 178.220 81.530 178.390 ;
        RECT 81.840 178.220 82.170 178.390 ;
        RECT 75.440 177.680 75.770 177.850 ;
        RECT 76.080 177.680 76.410 177.850 ;
        RECT 76.720 177.680 77.050 177.850 ;
        RECT 77.360 177.680 77.690 177.850 ;
        RECT 78.000 177.680 78.330 177.850 ;
        RECT 78.640 177.680 78.970 177.850 ;
        RECT 79.280 177.680 79.610 177.850 ;
        RECT 79.920 177.680 80.250 177.850 ;
        RECT 80.560 177.680 80.890 177.850 ;
        RECT 81.200 177.680 81.530 177.850 ;
        RECT 81.840 177.680 82.170 177.850 ;
        RECT 75.200 168.905 75.370 175.985 ;
        RECT 75.840 168.905 76.010 175.985 ;
        RECT 76.480 168.905 76.650 175.985 ;
        RECT 77.120 168.905 77.290 175.985 ;
        RECT 77.760 168.905 77.930 175.985 ;
        RECT 78.400 168.905 78.570 175.985 ;
        RECT 79.040 168.905 79.210 175.985 ;
        RECT 79.680 168.905 79.850 175.985 ;
        RECT 80.320 168.905 80.490 175.985 ;
        RECT 80.960 168.905 81.130 175.985 ;
        RECT 81.600 168.905 81.770 175.985 ;
        RECT 82.240 168.905 82.410 175.985 ;
        RECT 75.440 167.040 75.770 167.210 ;
        RECT 76.080 167.040 76.410 167.210 ;
        RECT 76.720 167.040 77.050 167.210 ;
        RECT 77.360 167.040 77.690 167.210 ;
        RECT 78.000 167.040 78.330 167.210 ;
        RECT 78.640 167.040 78.970 167.210 ;
        RECT 79.280 167.040 79.610 167.210 ;
        RECT 79.920 167.040 80.250 167.210 ;
        RECT 80.560 167.040 80.890 167.210 ;
        RECT 81.200 167.040 81.530 167.210 ;
        RECT 81.840 167.040 82.170 167.210 ;
        RECT 82.810 166.700 82.980 189.370 ;
        RECT 74.630 166.530 82.980 166.700 ;
        RECT 60.380 165.400 62.330 165.570 ;
        RECT 60.380 161.500 60.550 165.400 ;
        RECT 61.190 164.890 61.520 165.060 ;
        RECT 60.950 163.130 61.120 163.770 ;
        RECT 61.590 163.130 61.760 163.770 ;
        RECT 61.190 161.840 61.520 162.010 ;
        RECT 62.160 161.500 62.330 165.400 ;
        RECT 60.380 161.330 62.330 161.500 ;
        RECT 63.980 165.400 65.930 165.570 ;
        RECT 63.980 161.500 64.150 165.400 ;
        RECT 64.790 164.890 65.120 165.060 ;
        RECT 64.550 163.130 64.720 163.770 ;
        RECT 65.190 163.130 65.360 163.770 ;
        RECT 64.790 161.840 65.120 162.010 ;
        RECT 65.760 161.500 65.930 165.400 ;
        RECT 63.980 161.330 65.930 161.500 ;
        RECT 67.630 165.450 69.580 165.620 ;
        RECT 67.630 161.550 67.800 165.450 ;
        RECT 68.440 164.940 68.770 165.110 ;
        RECT 68.200 163.180 68.370 163.820 ;
        RECT 68.840 163.180 69.010 163.820 ;
        RECT 68.440 161.890 68.770 162.060 ;
        RECT 69.410 161.550 69.580 165.450 ;
        RECT 67.630 161.380 69.580 161.550 ;
        RECT 72.730 165.440 84.920 165.610 ;
        RECT 50.380 160.080 52.330 160.250 ;
        RECT 45.630 158.560 51.230 158.730 ;
        RECT 35.030 158.290 40.630 158.460 ;
        RECT 35.030 139.800 35.200 158.290 ;
        RECT 35.910 157.780 39.750 157.950 ;
        RECT 35.600 150.750 35.770 156.430 ;
        RECT 39.890 150.750 40.060 156.430 ;
        RECT 35.910 149.230 39.750 149.400 ;
        RECT 35.910 148.690 39.750 148.860 ;
        RECT 35.600 141.660 35.770 147.340 ;
        RECT 39.890 141.660 40.060 147.340 ;
        RECT 35.910 140.140 39.750 140.310 ;
        RECT 40.460 139.800 40.630 158.290 ;
        RECT 35.030 139.630 40.630 139.800 ;
        RECT 35.030 138.350 40.630 138.520 ;
        RECT 29.480 130.980 31.430 131.150 ;
        RECT 32.230 132.850 34.180 133.020 ;
        RECT 12.180 128.990 17.360 129.160 ;
        RECT 12.180 117.500 12.350 128.990 ;
        RECT 13.060 128.480 13.900 128.650 ;
        RECT 14.350 128.480 15.190 128.650 ;
        RECT 15.640 128.480 16.480 128.650 ;
        RECT 12.750 119.705 12.920 126.785 ;
        RECT 14.040 119.705 14.210 126.785 ;
        RECT 15.330 119.705 15.500 126.785 ;
        RECT 16.620 119.705 16.790 126.785 ;
        RECT 13.060 117.840 13.900 118.010 ;
        RECT 14.350 117.840 15.190 118.010 ;
        RECT 15.640 117.840 16.480 118.010 ;
        RECT 17.190 117.500 17.360 128.990 ;
        RECT 12.180 117.330 17.360 117.500 ;
        RECT 19.030 128.990 20.980 129.160 ;
        RECT 19.030 117.500 19.200 128.990 ;
        RECT 19.840 128.480 20.170 128.650 ;
        RECT 19.600 119.705 19.770 126.785 ;
        RECT 20.240 119.705 20.410 126.785 ;
        RECT 19.840 117.840 20.170 118.010 ;
        RECT 20.810 117.500 20.980 128.990 ;
        RECT 19.030 117.330 20.980 117.500 ;
        RECT 22.630 129.140 27.810 129.310 ;
        RECT 22.630 117.650 22.800 129.140 ;
        RECT 23.510 128.630 24.350 128.800 ;
        RECT 24.800 128.630 25.640 128.800 ;
        RECT 26.090 128.630 26.930 128.800 ;
        RECT 23.200 119.855 23.370 126.935 ;
        RECT 24.490 119.855 24.660 126.935 ;
        RECT 25.780 119.855 25.950 126.935 ;
        RECT 27.070 119.855 27.240 126.935 ;
        RECT 23.510 117.990 24.350 118.160 ;
        RECT 24.800 117.990 25.640 118.160 ;
        RECT 26.090 117.990 26.930 118.160 ;
        RECT 27.640 117.650 27.810 129.140 ;
        RECT 22.630 117.480 27.810 117.650 ;
        RECT 29.480 129.140 31.430 129.310 ;
        RECT 29.480 117.650 29.650 129.140 ;
        RECT 30.290 128.630 30.620 128.800 ;
        RECT 30.050 119.855 30.220 126.935 ;
        RECT 30.690 119.855 30.860 126.935 ;
        RECT 30.290 117.990 30.620 118.160 ;
        RECT 31.260 117.650 31.430 129.140 ;
        RECT 32.230 128.950 32.400 132.850 ;
        RECT 33.040 132.340 33.370 132.510 ;
        RECT 32.800 129.985 32.970 131.815 ;
        RECT 33.440 129.985 33.610 131.815 ;
        RECT 33.040 129.290 33.370 129.460 ;
        RECT 34.010 128.950 34.180 132.850 ;
        RECT 32.230 128.780 34.180 128.950 ;
        RECT 35.030 128.950 35.200 138.350 ;
        RECT 35.910 137.840 39.750 138.010 ;
        RECT 35.600 130.810 35.770 136.490 ;
        RECT 39.890 130.810 40.060 136.490 ;
        RECT 35.910 129.290 39.750 129.460 ;
        RECT 40.460 128.950 40.630 138.350 ;
        RECT 35.030 128.780 40.630 128.950 ;
        RECT 35.035 127.505 40.635 127.675 ;
        RECT 32.230 122.000 34.180 122.170 ;
        RECT 32.230 118.100 32.400 122.000 ;
        RECT 33.040 121.490 33.370 121.660 ;
        RECT 32.800 119.135 32.970 120.965 ;
        RECT 33.440 119.135 33.610 120.965 ;
        RECT 33.040 118.440 33.370 118.610 ;
        RECT 34.010 118.100 34.180 122.000 ;
        RECT 32.230 117.930 34.180 118.100 ;
        RECT 35.035 118.105 35.205 127.505 ;
        RECT 35.915 126.995 39.755 127.165 ;
        RECT 35.605 119.965 35.775 125.645 ;
        RECT 39.895 119.965 40.065 125.645 ;
        RECT 35.915 118.445 39.755 118.615 ;
        RECT 40.465 118.105 40.635 127.505 ;
        RECT 35.035 117.935 40.635 118.105 ;
        RECT 29.480 117.480 31.430 117.650 ;
        RECT 45.630 117.350 45.800 158.560 ;
        RECT 46.510 158.050 50.350 158.220 ;
        RECT 46.200 155.560 46.370 157.160 ;
        RECT 50.490 155.560 50.660 157.160 ;
        RECT 46.510 154.500 50.350 154.670 ;
        RECT 46.510 153.960 50.350 154.130 ;
        RECT 46.200 151.470 46.370 153.070 ;
        RECT 50.490 151.470 50.660 153.070 ;
        RECT 46.510 150.410 50.350 150.580 ;
        RECT 46.510 149.870 50.350 150.040 ;
        RECT 46.200 147.380 46.370 148.980 ;
        RECT 50.490 147.380 50.660 148.980 ;
        RECT 46.510 146.320 50.350 146.490 ;
        RECT 46.510 145.780 50.350 145.950 ;
        RECT 46.200 143.290 46.370 144.890 ;
        RECT 50.490 143.290 50.660 144.890 ;
        RECT 46.510 142.230 50.350 142.400 ;
        RECT 46.510 141.690 50.350 141.860 ;
        RECT 46.200 139.200 46.370 140.800 ;
        RECT 50.490 139.200 50.660 140.800 ;
        RECT 46.510 138.140 50.350 138.310 ;
        RECT 46.510 137.600 50.350 137.770 ;
        RECT 46.200 135.110 46.370 136.710 ;
        RECT 50.490 135.110 50.660 136.710 ;
        RECT 46.510 134.050 50.350 134.220 ;
        RECT 46.510 133.510 50.350 133.680 ;
        RECT 46.200 131.020 46.370 132.620 ;
        RECT 50.490 131.020 50.660 132.620 ;
        RECT 46.510 129.960 50.350 130.130 ;
        RECT 46.510 129.420 50.350 129.590 ;
        RECT 46.200 126.930 46.370 128.530 ;
        RECT 50.490 126.930 50.660 128.530 ;
        RECT 46.510 125.870 50.350 126.040 ;
        RECT 46.510 125.330 50.350 125.500 ;
        RECT 46.200 122.840 46.370 124.440 ;
        RECT 50.490 122.840 50.660 124.440 ;
        RECT 46.510 121.780 50.350 121.950 ;
        RECT 46.510 121.240 50.350 121.410 ;
        RECT 46.200 118.750 46.370 120.350 ;
        RECT 50.490 118.750 50.660 120.350 ;
        RECT 46.510 117.690 50.350 117.860 ;
        RECT 51.060 117.350 51.230 158.560 ;
        RECT 72.730 157.950 72.900 165.440 ;
        RECT 73.540 164.930 73.870 165.100 ;
        RECT 74.180 164.930 74.510 165.100 ;
        RECT 74.820 164.930 75.150 165.100 ;
        RECT 75.460 164.930 75.790 165.100 ;
        RECT 76.100 164.930 76.430 165.100 ;
        RECT 76.740 164.930 77.070 165.100 ;
        RECT 77.380 164.930 77.710 165.100 ;
        RECT 78.020 164.930 78.350 165.100 ;
        RECT 78.660 164.930 78.990 165.100 ;
        RECT 79.300 164.930 79.630 165.100 ;
        RECT 79.940 164.930 80.270 165.100 ;
        RECT 80.580 164.930 80.910 165.100 ;
        RECT 81.220 164.930 81.550 165.100 ;
        RECT 81.860 164.930 82.190 165.100 ;
        RECT 82.500 164.930 82.830 165.100 ;
        RECT 83.140 164.930 83.470 165.100 ;
        RECT 83.780 164.930 84.110 165.100 ;
        RECT 73.300 163.170 73.470 163.810 ;
        RECT 73.940 163.170 74.110 163.810 ;
        RECT 74.580 163.170 74.750 163.810 ;
        RECT 75.220 163.170 75.390 163.810 ;
        RECT 75.860 163.170 76.030 163.810 ;
        RECT 76.500 163.170 76.670 163.810 ;
        RECT 77.140 163.170 77.310 163.810 ;
        RECT 77.780 163.170 77.950 163.810 ;
        RECT 78.420 163.170 78.590 163.810 ;
        RECT 79.060 163.170 79.230 163.810 ;
        RECT 79.700 163.170 79.870 163.810 ;
        RECT 80.340 163.170 80.510 163.810 ;
        RECT 80.980 163.170 81.150 163.810 ;
        RECT 81.620 163.170 81.790 163.810 ;
        RECT 82.260 163.170 82.430 163.810 ;
        RECT 82.900 163.170 83.070 163.810 ;
        RECT 83.540 163.170 83.710 163.810 ;
        RECT 84.180 163.170 84.350 163.810 ;
        RECT 73.540 161.880 73.870 162.050 ;
        RECT 74.180 161.880 74.510 162.050 ;
        RECT 74.820 161.880 75.150 162.050 ;
        RECT 75.460 161.880 75.790 162.050 ;
        RECT 76.100 161.880 76.430 162.050 ;
        RECT 76.740 161.880 77.070 162.050 ;
        RECT 77.380 161.880 77.710 162.050 ;
        RECT 78.020 161.880 78.350 162.050 ;
        RECT 78.660 161.880 78.990 162.050 ;
        RECT 79.300 161.880 79.630 162.050 ;
        RECT 79.940 161.880 80.270 162.050 ;
        RECT 80.580 161.880 80.910 162.050 ;
        RECT 81.220 161.880 81.550 162.050 ;
        RECT 81.860 161.880 82.190 162.050 ;
        RECT 82.500 161.880 82.830 162.050 ;
        RECT 83.140 161.880 83.470 162.050 ;
        RECT 83.780 161.880 84.110 162.050 ;
        RECT 73.540 161.340 73.870 161.510 ;
        RECT 74.180 161.340 74.510 161.510 ;
        RECT 74.820 161.340 75.150 161.510 ;
        RECT 75.460 161.340 75.790 161.510 ;
        RECT 76.100 161.340 76.430 161.510 ;
        RECT 76.740 161.340 77.070 161.510 ;
        RECT 77.380 161.340 77.710 161.510 ;
        RECT 78.020 161.340 78.350 161.510 ;
        RECT 78.660 161.340 78.990 161.510 ;
        RECT 79.300 161.340 79.630 161.510 ;
        RECT 79.940 161.340 80.270 161.510 ;
        RECT 80.580 161.340 80.910 161.510 ;
        RECT 81.220 161.340 81.550 161.510 ;
        RECT 81.860 161.340 82.190 161.510 ;
        RECT 82.500 161.340 82.830 161.510 ;
        RECT 83.140 161.340 83.470 161.510 ;
        RECT 83.780 161.340 84.110 161.510 ;
        RECT 73.300 159.580 73.470 160.220 ;
        RECT 73.940 159.580 74.110 160.220 ;
        RECT 74.580 159.580 74.750 160.220 ;
        RECT 75.220 159.580 75.390 160.220 ;
        RECT 75.860 159.580 76.030 160.220 ;
        RECT 76.500 159.580 76.670 160.220 ;
        RECT 77.140 159.580 77.310 160.220 ;
        RECT 77.780 159.580 77.950 160.220 ;
        RECT 78.420 159.580 78.590 160.220 ;
        RECT 79.060 159.580 79.230 160.220 ;
        RECT 79.700 159.580 79.870 160.220 ;
        RECT 80.340 159.580 80.510 160.220 ;
        RECT 80.980 159.580 81.150 160.220 ;
        RECT 81.620 159.580 81.790 160.220 ;
        RECT 82.260 159.580 82.430 160.220 ;
        RECT 82.900 159.580 83.070 160.220 ;
        RECT 83.540 159.580 83.710 160.220 ;
        RECT 84.180 159.580 84.350 160.220 ;
        RECT 73.540 158.290 73.870 158.460 ;
        RECT 74.180 158.290 74.510 158.460 ;
        RECT 74.820 158.290 75.150 158.460 ;
        RECT 75.460 158.290 75.790 158.460 ;
        RECT 76.100 158.290 76.430 158.460 ;
        RECT 76.740 158.290 77.070 158.460 ;
        RECT 77.380 158.290 77.710 158.460 ;
        RECT 78.020 158.290 78.350 158.460 ;
        RECT 78.660 158.290 78.990 158.460 ;
        RECT 79.300 158.290 79.630 158.460 ;
        RECT 79.940 158.290 80.270 158.460 ;
        RECT 80.580 158.290 80.910 158.460 ;
        RECT 81.220 158.290 81.550 158.460 ;
        RECT 81.860 158.290 82.190 158.460 ;
        RECT 82.500 158.290 82.830 158.460 ;
        RECT 83.140 158.290 83.470 158.460 ;
        RECT 83.780 158.290 84.110 158.460 ;
        RECT 84.750 157.950 84.920 165.440 ;
        RECT 72.730 157.780 84.920 157.950 ;
        RECT 75.180 149.690 77.780 149.860 ;
        RECT 75.180 146.600 75.350 149.690 ;
        RECT 75.750 147.560 75.920 149.040 ;
        RECT 77.040 147.560 77.210 149.040 ;
        RECT 76.060 146.940 76.900 147.110 ;
        RECT 77.610 146.600 77.780 149.690 ;
        RECT 75.180 146.430 77.780 146.600 ;
        RECT 79.430 149.690 82.030 149.860 ;
        RECT 79.430 146.600 79.600 149.690 ;
        RECT 80.000 147.560 80.170 149.040 ;
        RECT 81.290 147.560 81.460 149.040 ;
        RECT 80.310 146.940 81.150 147.110 ;
        RECT 81.860 146.600 82.030 149.690 ;
        RECT 79.430 146.430 82.030 146.600 ;
        RECT 74.480 144.990 77.770 145.160 ;
        RECT 45.630 117.180 51.230 117.350 ;
        RECT 53.280 134.760 58.880 134.930 ;
        RECT 23.130 115.660 25.730 115.665 ;
        RECT 12.300 115.490 17.330 115.660 ;
        RECT 12.300 106.350 12.470 115.490 ;
        RECT 13.100 114.975 14.100 115.145 ;
        RECT 12.870 106.720 13.040 114.760 ;
        RECT 14.160 106.720 14.330 114.760 ;
        RECT 14.730 106.350 14.900 115.490 ;
        RECT 15.530 114.975 16.530 115.145 ;
        RECT 15.300 106.720 15.470 114.760 ;
        RECT 16.590 106.720 16.760 114.760 ;
        RECT 17.160 106.350 17.330 115.490 ;
        RECT 12.300 106.180 17.330 106.350 ;
        RECT 17.700 115.440 20.300 115.610 ;
        RECT 17.700 106.350 17.870 115.440 ;
        RECT 18.500 114.930 19.500 115.100 ;
        RECT 18.270 106.720 18.440 114.760 ;
        RECT 19.560 106.720 19.730 114.760 ;
        RECT 20.130 106.350 20.300 115.440 ;
        RECT 17.700 106.180 20.300 106.350 ;
        RECT 20.700 115.495 25.730 115.660 ;
        RECT 20.700 115.490 23.300 115.495 ;
        RECT 20.700 106.350 20.870 115.490 ;
        RECT 21.500 114.975 22.500 115.145 ;
        RECT 21.270 106.720 21.440 114.760 ;
        RECT 22.560 106.720 22.730 114.760 ;
        RECT 23.130 106.355 23.300 115.490 ;
        RECT 23.930 114.980 24.930 115.150 ;
        RECT 23.700 106.725 23.870 114.765 ;
        RECT 24.990 106.725 25.160 114.765 ;
        RECT 25.560 106.355 25.730 115.495 ;
        RECT 23.130 106.350 25.730 106.355 ;
        RECT 20.700 106.185 25.730 106.350 ;
        RECT 26.110 115.455 28.710 115.625 ;
        RECT 26.110 106.365 26.280 115.455 ;
        RECT 26.910 114.945 27.910 115.115 ;
        RECT 26.680 106.735 26.850 114.775 ;
        RECT 27.970 106.735 28.140 114.775 ;
        RECT 28.540 106.365 28.710 115.455 ;
        RECT 26.110 106.195 28.710 106.365 ;
        RECT 29.100 115.490 38.895 115.660 ;
        RECT 29.100 106.350 29.270 115.490 ;
        RECT 29.900 114.975 30.900 115.145 ;
        RECT 29.670 106.720 29.840 114.760 ;
        RECT 30.960 106.720 31.130 114.760 ;
        RECT 31.500 106.350 31.700 115.490 ;
        RECT 32.300 114.975 33.300 115.145 ;
        RECT 32.070 106.720 32.240 114.760 ;
        RECT 33.360 106.720 33.530 114.760 ;
        RECT 33.900 106.350 34.100 115.490 ;
        RECT 34.700 114.975 35.700 115.145 ;
        RECT 34.470 106.720 34.640 114.760 ;
        RECT 35.760 106.720 35.930 114.760 ;
        RECT 36.295 106.350 36.500 115.490 ;
        RECT 37.095 114.975 38.095 115.145 ;
        RECT 36.865 106.720 37.035 114.760 ;
        RECT 38.155 106.720 38.325 114.760 ;
        RECT 38.725 111.080 38.895 115.490 ;
        RECT 39.300 113.160 48.900 113.330 ;
        RECT 39.300 111.650 39.470 113.160 ;
        RECT 40.100 112.650 48.100 112.820 ;
        RECT 39.870 112.020 40.040 112.480 ;
        RECT 48.160 112.020 48.330 112.480 ;
        RECT 48.730 111.650 48.900 113.160 ;
        RECT 39.300 111.480 48.900 111.650 ;
        RECT 38.725 110.910 48.400 111.080 ;
        RECT 38.725 109.350 38.970 110.910 ;
        RECT 39.600 110.395 47.600 110.565 ;
        RECT 39.370 109.720 39.540 110.180 ;
        RECT 47.660 109.720 47.830 110.180 ;
        RECT 48.230 109.350 48.400 110.910 ;
        RECT 38.725 109.180 48.400 109.350 ;
        RECT 38.725 106.350 38.895 109.180 ;
        RECT 20.700 106.180 23.300 106.185 ;
        RECT 29.100 106.180 38.895 106.350 ;
        RECT 39.300 108.610 48.730 108.780 ;
        RECT 39.300 106.350 39.470 108.610 ;
        RECT 39.840 108.040 47.880 108.210 ;
        RECT 48.050 106.980 48.220 107.980 ;
        RECT 39.840 106.750 47.880 106.920 ;
        RECT 48.560 106.350 48.730 108.610 ;
        RECT 39.300 106.180 48.730 106.350 ;
        RECT 12.280 105.410 34.320 105.510 ;
        RECT 12.280 105.340 48.900 105.410 ;
        RECT 12.280 96.250 12.450 105.340 ;
        RECT 13.080 104.830 14.080 105.000 ;
        RECT 12.850 96.620 13.020 104.660 ;
        RECT 14.140 96.620 14.310 104.660 ;
        RECT 14.710 96.250 14.880 105.340 ;
        RECT 15.510 104.830 16.510 105.000 ;
        RECT 15.280 96.620 15.450 104.660 ;
        RECT 16.570 96.620 16.740 104.660 ;
        RECT 17.140 96.250 17.310 105.340 ;
        RECT 17.940 104.830 18.940 105.000 ;
        RECT 17.710 96.620 17.880 104.660 ;
        RECT 19.000 96.620 19.170 104.660 ;
        RECT 19.570 96.250 19.740 105.340 ;
        RECT 20.370 104.830 21.370 105.000 ;
        RECT 20.140 96.620 20.310 104.660 ;
        RECT 21.430 96.620 21.600 104.660 ;
        RECT 22.000 96.250 22.170 105.340 ;
        RECT 22.800 104.830 23.800 105.000 ;
        RECT 22.570 96.620 22.740 104.660 ;
        RECT 23.860 96.620 24.030 104.660 ;
        RECT 24.430 96.250 24.600 105.340 ;
        RECT 25.230 104.830 26.230 105.000 ;
        RECT 25.000 96.620 25.170 104.660 ;
        RECT 26.290 96.620 26.460 104.660 ;
        RECT 26.860 96.250 27.030 105.340 ;
        RECT 27.660 104.830 28.660 105.000 ;
        RECT 27.430 96.620 27.600 104.660 ;
        RECT 28.720 96.620 28.890 104.660 ;
        RECT 29.290 96.250 29.460 105.340 ;
        RECT 30.090 104.830 31.090 105.000 ;
        RECT 29.860 96.620 30.030 104.660 ;
        RECT 31.150 96.620 31.320 104.660 ;
        RECT 31.720 96.250 31.890 105.340 ;
        RECT 34.150 105.240 48.900 105.340 ;
        RECT 32.520 104.830 33.520 105.000 ;
        RECT 32.290 96.620 32.460 104.660 ;
        RECT 33.580 96.620 33.750 104.660 ;
        RECT 34.150 103.150 34.370 105.240 ;
        RECT 35.000 104.730 48.100 104.900 ;
        RECT 34.770 103.520 34.940 104.560 ;
        RECT 48.160 103.520 48.330 104.560 ;
        RECT 48.730 103.150 48.900 105.240 ;
        RECT 34.150 102.980 48.900 103.150 ;
        RECT 34.150 102.940 43.800 102.980 ;
        RECT 34.150 100.850 34.370 102.940 ;
        RECT 35.000 102.430 43.000 102.600 ;
        RECT 34.770 101.220 34.940 102.260 ;
        RECT 43.060 101.220 43.230 102.260 ;
        RECT 43.630 100.850 43.800 102.940 ;
        RECT 34.150 100.640 43.800 100.850 ;
        RECT 34.150 98.550 34.370 100.640 ;
        RECT 35.000 100.130 43.000 100.300 ;
        RECT 34.770 98.920 34.940 99.960 ;
        RECT 43.060 98.920 43.230 99.960 ;
        RECT 43.630 98.550 43.800 100.640 ;
        RECT 34.150 98.340 43.800 98.550 ;
        RECT 34.150 96.250 34.370 98.340 ;
        RECT 35.000 97.830 43.000 98.000 ;
        RECT 34.770 96.620 34.940 97.660 ;
        RECT 43.060 96.620 43.230 97.660 ;
        RECT 43.630 96.250 43.800 98.340 ;
        RECT 12.280 96.080 43.800 96.250 ;
        RECT 53.280 93.550 53.450 134.760 ;
        RECT 54.160 134.250 58.000 134.420 ;
        RECT 53.850 131.760 54.020 133.360 ;
        RECT 58.140 131.760 58.310 133.360 ;
        RECT 54.160 130.700 58.000 130.870 ;
        RECT 54.160 130.160 58.000 130.330 ;
        RECT 53.850 127.670 54.020 129.270 ;
        RECT 58.140 127.670 58.310 129.270 ;
        RECT 54.160 126.610 58.000 126.780 ;
        RECT 54.160 126.070 58.000 126.240 ;
        RECT 53.850 123.580 54.020 125.180 ;
        RECT 58.140 123.580 58.310 125.180 ;
        RECT 54.160 122.520 58.000 122.690 ;
        RECT 54.160 121.980 58.000 122.150 ;
        RECT 53.850 119.490 54.020 121.090 ;
        RECT 58.140 119.490 58.310 121.090 ;
        RECT 54.160 118.430 58.000 118.600 ;
        RECT 54.160 117.890 58.000 118.060 ;
        RECT 53.850 115.400 54.020 117.000 ;
        RECT 58.140 115.400 58.310 117.000 ;
        RECT 54.160 114.340 58.000 114.510 ;
        RECT 54.160 113.800 58.000 113.970 ;
        RECT 53.850 111.310 54.020 112.910 ;
        RECT 58.140 111.310 58.310 112.910 ;
        RECT 54.160 110.250 58.000 110.420 ;
        RECT 54.160 109.710 58.000 109.880 ;
        RECT 53.850 107.220 54.020 108.820 ;
        RECT 58.140 107.220 58.310 108.820 ;
        RECT 54.160 106.160 58.000 106.330 ;
        RECT 54.160 105.620 58.000 105.790 ;
        RECT 53.850 103.130 54.020 104.730 ;
        RECT 58.140 103.130 58.310 104.730 ;
        RECT 54.160 102.070 58.000 102.240 ;
        RECT 54.160 101.530 58.000 101.700 ;
        RECT 53.850 99.040 54.020 100.640 ;
        RECT 58.140 99.040 58.310 100.640 ;
        RECT 54.160 97.980 58.000 98.150 ;
        RECT 54.160 97.440 58.000 97.610 ;
        RECT 53.850 94.950 54.020 96.550 ;
        RECT 58.140 94.950 58.310 96.550 ;
        RECT 54.160 93.890 58.000 94.060 ;
        RECT 58.710 93.550 58.880 134.760 ;
        RECT 74.480 133.500 74.650 144.990 ;
        RECT 75.360 144.480 75.900 144.650 ;
        RECT 76.350 144.480 76.890 144.650 ;
        RECT 75.050 135.705 75.220 142.785 ;
        RECT 76.040 135.705 76.210 142.785 ;
        RECT 77.030 135.705 77.200 142.785 ;
        RECT 75.360 133.840 75.900 134.010 ;
        RECT 76.350 133.840 76.890 134.010 ;
        RECT 77.600 133.500 77.770 144.990 ;
        RECT 74.480 133.330 77.770 133.500 ;
        RECT 79.430 144.990 82.720 145.160 ;
        RECT 79.430 133.500 79.600 144.990 ;
        RECT 80.310 144.480 80.850 144.650 ;
        RECT 81.300 144.480 81.840 144.650 ;
        RECT 80.000 135.705 80.170 142.785 ;
        RECT 80.990 135.705 81.160 142.785 ;
        RECT 81.980 135.705 82.150 142.785 ;
        RECT 80.310 133.840 80.850 134.010 ;
        RECT 81.300 133.840 81.840 134.010 ;
        RECT 82.550 133.500 82.720 144.990 ;
        RECT 79.430 133.330 82.720 133.500 ;
        RECT 59.880 131.600 77.770 131.770 ;
        RECT 59.880 110.200 60.050 131.600 ;
        RECT 60.760 131.090 68.600 131.260 ;
        RECT 69.050 131.090 76.890 131.260 ;
        RECT 60.450 113.860 60.620 127.940 ;
        RECT 68.740 113.860 68.910 127.940 ;
        RECT 77.030 113.860 77.200 127.940 ;
        RECT 60.760 110.540 68.600 110.710 ;
        RECT 69.050 110.540 76.890 110.710 ;
        RECT 77.600 110.200 77.770 131.600 ;
        RECT 59.880 110.030 77.770 110.200 ;
        RECT 79.430 131.600 97.320 131.770 ;
        RECT 79.430 110.200 79.600 131.600 ;
        RECT 80.310 131.090 88.150 131.260 ;
        RECT 88.600 131.090 96.440 131.260 ;
        RECT 80.000 113.860 80.170 127.940 ;
        RECT 88.290 113.860 88.460 127.940 ;
        RECT 96.580 113.860 96.750 127.940 ;
        RECT 80.310 110.540 88.150 110.710 ;
        RECT 88.600 110.540 96.440 110.710 ;
        RECT 97.150 110.200 97.320 131.600 ;
        RECT 98.430 129.940 100.380 130.110 ;
        RECT 98.430 118.450 98.600 129.940 ;
        RECT 99.240 129.430 99.570 129.600 ;
        RECT 99.000 120.655 99.170 127.735 ;
        RECT 99.640 120.655 99.810 127.735 ;
        RECT 99.240 118.790 99.570 118.960 ;
        RECT 100.210 118.450 100.380 129.940 ;
        RECT 98.430 118.280 100.380 118.450 ;
        RECT 102.030 129.940 103.980 130.110 ;
        RECT 102.030 118.450 102.200 129.940 ;
        RECT 102.840 129.430 103.170 129.600 ;
        RECT 102.600 120.655 102.770 127.735 ;
        RECT 103.240 120.655 103.410 127.735 ;
        RECT 102.840 118.790 103.170 118.960 ;
        RECT 103.810 118.450 103.980 129.940 ;
        RECT 102.030 118.280 103.980 118.450 ;
        RECT 105.630 129.940 107.580 130.110 ;
        RECT 105.630 118.450 105.800 129.940 ;
        RECT 106.440 129.430 106.770 129.600 ;
        RECT 106.200 120.655 106.370 127.735 ;
        RECT 106.840 120.655 107.010 127.735 ;
        RECT 106.440 118.790 106.770 118.960 ;
        RECT 107.410 118.450 107.580 129.940 ;
        RECT 105.630 118.280 107.580 118.450 ;
        RECT 109.230 122.440 111.180 122.610 ;
        RECT 109.230 118.450 109.400 122.440 ;
        RECT 110.040 121.930 110.370 122.100 ;
        RECT 109.800 119.530 109.970 121.360 ;
        RECT 110.440 119.530 110.610 121.360 ;
        RECT 110.040 118.790 110.370 118.960 ;
        RECT 111.010 118.450 111.180 122.440 ;
        RECT 109.230 118.280 111.180 118.450 ;
        RECT 79.430 110.030 97.320 110.200 ;
        RECT 98.430 117.250 116.320 117.420 ;
        RECT 53.280 93.380 58.880 93.550 ;
        RECT 59.880 108.200 77.770 108.370 ;
        RECT 46.880 90.200 52.480 90.370 ;
        RECT 46.880 85.800 47.050 90.200 ;
        RECT 47.760 89.690 51.600 89.860 ;
        RECT 47.450 87.200 47.620 88.800 ;
        RECT 51.740 87.200 51.910 88.800 ;
        RECT 47.760 86.140 51.600 86.310 ;
        RECT 52.310 85.800 52.480 90.200 ;
        RECT 46.880 85.630 52.480 85.800 ;
        RECT 53.280 90.200 58.880 90.370 ;
        RECT 53.280 85.800 53.450 90.200 ;
        RECT 54.160 89.690 58.000 89.860 ;
        RECT 53.850 87.200 54.020 88.800 ;
        RECT 58.140 87.200 58.310 88.800 ;
        RECT 54.160 86.140 58.000 86.310 ;
        RECT 58.710 85.800 58.880 90.200 ;
        RECT 59.880 86.800 60.050 108.200 ;
        RECT 60.760 107.690 68.600 107.860 ;
        RECT 69.050 107.690 76.890 107.860 ;
        RECT 60.450 90.460 60.620 104.540 ;
        RECT 68.740 90.460 68.910 104.540 ;
        RECT 77.030 90.460 77.200 104.540 ;
        RECT 60.760 87.140 68.600 87.310 ;
        RECT 69.050 87.140 76.890 87.310 ;
        RECT 77.600 86.800 77.770 108.200 ;
        RECT 59.880 86.630 77.770 86.800 ;
        RECT 79.430 108.200 97.320 108.370 ;
        RECT 79.430 86.800 79.600 108.200 ;
        RECT 80.310 107.690 88.150 107.860 ;
        RECT 88.600 107.690 96.440 107.860 ;
        RECT 80.000 90.460 80.170 104.540 ;
        RECT 88.290 90.460 88.460 104.540 ;
        RECT 96.580 90.460 96.750 104.540 ;
        RECT 80.310 87.140 88.150 87.310 ;
        RECT 88.600 87.140 96.440 87.310 ;
        RECT 97.150 86.800 97.320 108.200 ;
        RECT 98.430 95.850 98.600 117.250 ;
        RECT 99.310 116.740 107.150 116.910 ;
        RECT 107.600 116.740 115.440 116.910 ;
        RECT 99.000 99.510 99.170 113.590 ;
        RECT 107.290 99.510 107.460 113.590 ;
        RECT 115.580 99.510 115.750 113.590 ;
        RECT 99.310 96.190 107.150 96.360 ;
        RECT 107.600 96.190 115.440 96.360 ;
        RECT 116.150 95.850 116.320 117.250 ;
        RECT 98.430 95.680 116.320 95.850 ;
        RECT 79.430 86.630 97.320 86.800 ;
        RECT 53.280 85.630 58.880 85.800 ;
        RECT 44.780 84.790 77.770 84.960 ;
        RECT 44.780 63.300 44.950 84.790 ;
        RECT 45.660 84.280 46.200 84.450 ;
        RECT 46.650 84.280 47.190 84.450 ;
        RECT 47.640 84.280 48.180 84.450 ;
        RECT 48.630 84.280 49.170 84.450 ;
        RECT 49.620 84.280 50.160 84.450 ;
        RECT 50.610 84.280 51.150 84.450 ;
        RECT 51.600 84.280 52.140 84.450 ;
        RECT 52.590 84.280 53.130 84.450 ;
        RECT 53.580 84.280 54.120 84.450 ;
        RECT 54.570 84.280 55.110 84.450 ;
        RECT 55.560 84.280 56.100 84.450 ;
        RECT 56.550 84.280 57.090 84.450 ;
        RECT 57.540 84.280 58.080 84.450 ;
        RECT 58.530 84.280 59.070 84.450 ;
        RECT 59.520 84.280 60.060 84.450 ;
        RECT 60.510 84.280 61.050 84.450 ;
        RECT 61.500 84.280 62.040 84.450 ;
        RECT 62.490 84.280 63.030 84.450 ;
        RECT 63.480 84.280 64.020 84.450 ;
        RECT 64.470 84.280 65.010 84.450 ;
        RECT 65.460 84.280 66.000 84.450 ;
        RECT 66.450 84.280 66.990 84.450 ;
        RECT 67.440 84.280 67.980 84.450 ;
        RECT 68.430 84.280 68.970 84.450 ;
        RECT 69.420 84.280 69.960 84.450 ;
        RECT 70.410 84.280 70.950 84.450 ;
        RECT 71.400 84.280 71.940 84.450 ;
        RECT 72.390 84.280 72.930 84.450 ;
        RECT 73.380 84.280 73.920 84.450 ;
        RECT 74.370 84.280 74.910 84.450 ;
        RECT 75.360 84.280 75.900 84.450 ;
        RECT 76.350 84.280 76.890 84.450 ;
        RECT 45.350 67.005 45.520 81.085 ;
        RECT 46.340 67.005 46.510 81.085 ;
        RECT 47.330 67.005 47.500 81.085 ;
        RECT 48.320 67.005 48.490 81.085 ;
        RECT 49.310 67.005 49.480 81.085 ;
        RECT 50.300 67.005 50.470 81.085 ;
        RECT 51.290 67.005 51.460 81.085 ;
        RECT 52.280 67.005 52.450 81.085 ;
        RECT 53.270 67.005 53.440 81.085 ;
        RECT 54.260 67.005 54.430 81.085 ;
        RECT 55.250 67.005 55.420 81.085 ;
        RECT 56.240 67.005 56.410 81.085 ;
        RECT 57.230 67.005 57.400 81.085 ;
        RECT 58.220 67.005 58.390 81.085 ;
        RECT 59.210 67.005 59.380 81.085 ;
        RECT 60.200 67.005 60.370 81.085 ;
        RECT 61.190 67.005 61.360 81.085 ;
        RECT 62.180 67.005 62.350 81.085 ;
        RECT 63.170 67.005 63.340 81.085 ;
        RECT 64.160 67.005 64.330 81.085 ;
        RECT 65.150 67.005 65.320 81.085 ;
        RECT 66.140 67.005 66.310 81.085 ;
        RECT 67.130 67.005 67.300 81.085 ;
        RECT 68.120 67.005 68.290 81.085 ;
        RECT 69.110 67.005 69.280 81.085 ;
        RECT 70.100 67.005 70.270 81.085 ;
        RECT 71.090 67.005 71.260 81.085 ;
        RECT 72.080 67.005 72.250 81.085 ;
        RECT 73.070 67.005 73.240 81.085 ;
        RECT 74.060 67.005 74.230 81.085 ;
        RECT 75.050 67.005 75.220 81.085 ;
        RECT 76.040 67.005 76.210 81.085 ;
        RECT 77.030 67.005 77.200 81.085 ;
        RECT 45.660 63.640 46.200 63.810 ;
        RECT 46.650 63.640 47.190 63.810 ;
        RECT 47.640 63.640 48.180 63.810 ;
        RECT 48.630 63.640 49.170 63.810 ;
        RECT 49.620 63.640 50.160 63.810 ;
        RECT 50.610 63.640 51.150 63.810 ;
        RECT 51.600 63.640 52.140 63.810 ;
        RECT 52.590 63.640 53.130 63.810 ;
        RECT 53.580 63.640 54.120 63.810 ;
        RECT 54.570 63.640 55.110 63.810 ;
        RECT 55.560 63.640 56.100 63.810 ;
        RECT 56.550 63.640 57.090 63.810 ;
        RECT 57.540 63.640 58.080 63.810 ;
        RECT 58.530 63.640 59.070 63.810 ;
        RECT 59.520 63.640 60.060 63.810 ;
        RECT 60.510 63.640 61.050 63.810 ;
        RECT 61.500 63.640 62.040 63.810 ;
        RECT 62.490 63.640 63.030 63.810 ;
        RECT 63.480 63.640 64.020 63.810 ;
        RECT 64.470 63.640 65.010 63.810 ;
        RECT 65.460 63.640 66.000 63.810 ;
        RECT 66.450 63.640 66.990 63.810 ;
        RECT 67.440 63.640 67.980 63.810 ;
        RECT 68.430 63.640 68.970 63.810 ;
        RECT 69.420 63.640 69.960 63.810 ;
        RECT 70.410 63.640 70.950 63.810 ;
        RECT 71.400 63.640 71.940 63.810 ;
        RECT 72.390 63.640 72.930 63.810 ;
        RECT 73.380 63.640 73.920 63.810 ;
        RECT 74.370 63.640 74.910 63.810 ;
        RECT 75.360 63.640 75.900 63.810 ;
        RECT 76.350 63.640 76.890 63.810 ;
        RECT 77.600 63.300 77.770 84.790 ;
        RECT 44.780 63.130 77.770 63.300 ;
        RECT 79.430 84.790 112.420 84.960 ;
        RECT 79.430 63.300 79.600 84.790 ;
        RECT 80.310 84.280 80.850 84.450 ;
        RECT 81.300 84.280 81.840 84.450 ;
        RECT 82.290 84.280 82.830 84.450 ;
        RECT 83.280 84.280 83.820 84.450 ;
        RECT 84.270 84.280 84.810 84.450 ;
        RECT 85.260 84.280 85.800 84.450 ;
        RECT 86.250 84.280 86.790 84.450 ;
        RECT 87.240 84.280 87.780 84.450 ;
        RECT 88.230 84.280 88.770 84.450 ;
        RECT 89.220 84.280 89.760 84.450 ;
        RECT 90.210 84.280 90.750 84.450 ;
        RECT 91.200 84.280 91.740 84.450 ;
        RECT 92.190 84.280 92.730 84.450 ;
        RECT 93.180 84.280 93.720 84.450 ;
        RECT 94.170 84.280 94.710 84.450 ;
        RECT 95.160 84.280 95.700 84.450 ;
        RECT 96.150 84.280 96.690 84.450 ;
        RECT 97.140 84.280 97.680 84.450 ;
        RECT 98.130 84.280 98.670 84.450 ;
        RECT 99.120 84.280 99.660 84.450 ;
        RECT 100.110 84.280 100.650 84.450 ;
        RECT 101.100 84.280 101.640 84.450 ;
        RECT 102.090 84.280 102.630 84.450 ;
        RECT 103.080 84.280 103.620 84.450 ;
        RECT 104.070 84.280 104.610 84.450 ;
        RECT 105.060 84.280 105.600 84.450 ;
        RECT 106.050 84.280 106.590 84.450 ;
        RECT 107.040 84.280 107.580 84.450 ;
        RECT 108.030 84.280 108.570 84.450 ;
        RECT 109.020 84.280 109.560 84.450 ;
        RECT 110.010 84.280 110.550 84.450 ;
        RECT 111.000 84.280 111.540 84.450 ;
        RECT 80.000 67.005 80.170 81.085 ;
        RECT 80.990 67.005 81.160 81.085 ;
        RECT 81.980 67.005 82.150 81.085 ;
        RECT 82.970 67.005 83.140 81.085 ;
        RECT 83.960 67.005 84.130 81.085 ;
        RECT 84.950 67.005 85.120 81.085 ;
        RECT 85.940 67.005 86.110 81.085 ;
        RECT 86.930 67.005 87.100 81.085 ;
        RECT 87.920 67.005 88.090 81.085 ;
        RECT 88.910 67.005 89.080 81.085 ;
        RECT 89.900 67.005 90.070 81.085 ;
        RECT 90.890 67.005 91.060 81.085 ;
        RECT 91.880 67.005 92.050 81.085 ;
        RECT 92.870 67.005 93.040 81.085 ;
        RECT 93.860 67.005 94.030 81.085 ;
        RECT 94.850 67.005 95.020 81.085 ;
        RECT 95.840 67.005 96.010 81.085 ;
        RECT 96.830 67.005 97.000 81.085 ;
        RECT 97.820 67.005 97.990 81.085 ;
        RECT 98.810 67.005 98.980 81.085 ;
        RECT 99.800 67.005 99.970 81.085 ;
        RECT 100.790 67.005 100.960 81.085 ;
        RECT 101.780 67.005 101.950 81.085 ;
        RECT 102.770 67.005 102.940 81.085 ;
        RECT 103.760 67.005 103.930 81.085 ;
        RECT 104.750 67.005 104.920 81.085 ;
        RECT 105.740 67.005 105.910 81.085 ;
        RECT 106.730 67.005 106.900 81.085 ;
        RECT 107.720 67.005 107.890 81.085 ;
        RECT 108.710 67.005 108.880 81.085 ;
        RECT 109.700 67.005 109.870 81.085 ;
        RECT 110.690 67.005 110.860 81.085 ;
        RECT 111.680 67.005 111.850 81.085 ;
        RECT 80.310 63.640 80.850 63.810 ;
        RECT 81.300 63.640 81.840 63.810 ;
        RECT 82.290 63.640 82.830 63.810 ;
        RECT 83.280 63.640 83.820 63.810 ;
        RECT 84.270 63.640 84.810 63.810 ;
        RECT 85.260 63.640 85.800 63.810 ;
        RECT 86.250 63.640 86.790 63.810 ;
        RECT 87.240 63.640 87.780 63.810 ;
        RECT 88.230 63.640 88.770 63.810 ;
        RECT 89.220 63.640 89.760 63.810 ;
        RECT 90.210 63.640 90.750 63.810 ;
        RECT 91.200 63.640 91.740 63.810 ;
        RECT 92.190 63.640 92.730 63.810 ;
        RECT 93.180 63.640 93.720 63.810 ;
        RECT 94.170 63.640 94.710 63.810 ;
        RECT 95.160 63.640 95.700 63.810 ;
        RECT 96.150 63.640 96.690 63.810 ;
        RECT 97.140 63.640 97.680 63.810 ;
        RECT 98.130 63.640 98.670 63.810 ;
        RECT 99.120 63.640 99.660 63.810 ;
        RECT 100.110 63.640 100.650 63.810 ;
        RECT 101.100 63.640 101.640 63.810 ;
        RECT 102.090 63.640 102.630 63.810 ;
        RECT 103.080 63.640 103.620 63.810 ;
        RECT 104.070 63.640 104.610 63.810 ;
        RECT 105.060 63.640 105.600 63.810 ;
        RECT 106.050 63.640 106.590 63.810 ;
        RECT 107.040 63.640 107.580 63.810 ;
        RECT 108.030 63.640 108.570 63.810 ;
        RECT 109.020 63.640 109.560 63.810 ;
        RECT 110.010 63.640 110.550 63.810 ;
        RECT 111.000 63.640 111.540 63.810 ;
        RECT 112.250 63.300 112.420 84.790 ;
        RECT 79.430 63.130 112.420 63.300 ;
        RECT 44.780 61.290 77.770 61.460 ;
        RECT 44.780 39.800 44.950 61.290 ;
        RECT 45.660 60.780 46.200 60.950 ;
        RECT 46.650 60.780 47.190 60.950 ;
        RECT 47.640 60.780 48.180 60.950 ;
        RECT 48.630 60.780 49.170 60.950 ;
        RECT 49.620 60.780 50.160 60.950 ;
        RECT 50.610 60.780 51.150 60.950 ;
        RECT 51.600 60.780 52.140 60.950 ;
        RECT 52.590 60.780 53.130 60.950 ;
        RECT 53.580 60.780 54.120 60.950 ;
        RECT 54.570 60.780 55.110 60.950 ;
        RECT 55.560 60.780 56.100 60.950 ;
        RECT 56.550 60.780 57.090 60.950 ;
        RECT 57.540 60.780 58.080 60.950 ;
        RECT 58.530 60.780 59.070 60.950 ;
        RECT 59.520 60.780 60.060 60.950 ;
        RECT 60.510 60.780 61.050 60.950 ;
        RECT 61.500 60.780 62.040 60.950 ;
        RECT 62.490 60.780 63.030 60.950 ;
        RECT 63.480 60.780 64.020 60.950 ;
        RECT 64.470 60.780 65.010 60.950 ;
        RECT 65.460 60.780 66.000 60.950 ;
        RECT 66.450 60.780 66.990 60.950 ;
        RECT 67.440 60.780 67.980 60.950 ;
        RECT 68.430 60.780 68.970 60.950 ;
        RECT 69.420 60.780 69.960 60.950 ;
        RECT 70.410 60.780 70.950 60.950 ;
        RECT 71.400 60.780 71.940 60.950 ;
        RECT 72.390 60.780 72.930 60.950 ;
        RECT 73.380 60.780 73.920 60.950 ;
        RECT 74.370 60.780 74.910 60.950 ;
        RECT 75.360 60.780 75.900 60.950 ;
        RECT 76.350 60.780 76.890 60.950 ;
        RECT 45.350 43.505 45.520 57.585 ;
        RECT 46.340 43.505 46.510 57.585 ;
        RECT 47.330 43.505 47.500 57.585 ;
        RECT 48.320 43.505 48.490 57.585 ;
        RECT 49.310 43.505 49.480 57.585 ;
        RECT 50.300 43.505 50.470 57.585 ;
        RECT 51.290 43.505 51.460 57.585 ;
        RECT 52.280 43.505 52.450 57.585 ;
        RECT 53.270 43.505 53.440 57.585 ;
        RECT 54.260 43.505 54.430 57.585 ;
        RECT 55.250 43.505 55.420 57.585 ;
        RECT 56.240 43.505 56.410 57.585 ;
        RECT 57.230 43.505 57.400 57.585 ;
        RECT 58.220 43.505 58.390 57.585 ;
        RECT 59.210 43.505 59.380 57.585 ;
        RECT 60.200 43.505 60.370 57.585 ;
        RECT 61.190 43.505 61.360 57.585 ;
        RECT 62.180 43.505 62.350 57.585 ;
        RECT 63.170 43.505 63.340 57.585 ;
        RECT 64.160 43.505 64.330 57.585 ;
        RECT 65.150 43.505 65.320 57.585 ;
        RECT 66.140 43.505 66.310 57.585 ;
        RECT 67.130 43.505 67.300 57.585 ;
        RECT 68.120 43.505 68.290 57.585 ;
        RECT 69.110 43.505 69.280 57.585 ;
        RECT 70.100 43.505 70.270 57.585 ;
        RECT 71.090 43.505 71.260 57.585 ;
        RECT 72.080 43.505 72.250 57.585 ;
        RECT 73.070 43.505 73.240 57.585 ;
        RECT 74.060 43.505 74.230 57.585 ;
        RECT 75.050 43.505 75.220 57.585 ;
        RECT 76.040 43.505 76.210 57.585 ;
        RECT 77.030 43.505 77.200 57.585 ;
        RECT 45.660 40.140 46.200 40.310 ;
        RECT 46.650 40.140 47.190 40.310 ;
        RECT 47.640 40.140 48.180 40.310 ;
        RECT 48.630 40.140 49.170 40.310 ;
        RECT 49.620 40.140 50.160 40.310 ;
        RECT 50.610 40.140 51.150 40.310 ;
        RECT 51.600 40.140 52.140 40.310 ;
        RECT 52.590 40.140 53.130 40.310 ;
        RECT 53.580 40.140 54.120 40.310 ;
        RECT 54.570 40.140 55.110 40.310 ;
        RECT 55.560 40.140 56.100 40.310 ;
        RECT 56.550 40.140 57.090 40.310 ;
        RECT 57.540 40.140 58.080 40.310 ;
        RECT 58.530 40.140 59.070 40.310 ;
        RECT 59.520 40.140 60.060 40.310 ;
        RECT 60.510 40.140 61.050 40.310 ;
        RECT 61.500 40.140 62.040 40.310 ;
        RECT 62.490 40.140 63.030 40.310 ;
        RECT 63.480 40.140 64.020 40.310 ;
        RECT 64.470 40.140 65.010 40.310 ;
        RECT 65.460 40.140 66.000 40.310 ;
        RECT 66.450 40.140 66.990 40.310 ;
        RECT 67.440 40.140 67.980 40.310 ;
        RECT 68.430 40.140 68.970 40.310 ;
        RECT 69.420 40.140 69.960 40.310 ;
        RECT 70.410 40.140 70.950 40.310 ;
        RECT 71.400 40.140 71.940 40.310 ;
        RECT 72.390 40.140 72.930 40.310 ;
        RECT 73.380 40.140 73.920 40.310 ;
        RECT 74.370 40.140 74.910 40.310 ;
        RECT 75.360 40.140 75.900 40.310 ;
        RECT 76.350 40.140 76.890 40.310 ;
        RECT 77.600 39.800 77.770 61.290 ;
        RECT 44.780 39.630 77.770 39.800 ;
        RECT 79.430 61.290 112.420 61.460 ;
        RECT 79.430 39.800 79.600 61.290 ;
        RECT 80.310 60.780 80.850 60.950 ;
        RECT 81.300 60.780 81.840 60.950 ;
        RECT 82.290 60.780 82.830 60.950 ;
        RECT 83.280 60.780 83.820 60.950 ;
        RECT 84.270 60.780 84.810 60.950 ;
        RECT 85.260 60.780 85.800 60.950 ;
        RECT 86.250 60.780 86.790 60.950 ;
        RECT 87.240 60.780 87.780 60.950 ;
        RECT 88.230 60.780 88.770 60.950 ;
        RECT 89.220 60.780 89.760 60.950 ;
        RECT 90.210 60.780 90.750 60.950 ;
        RECT 91.200 60.780 91.740 60.950 ;
        RECT 92.190 60.780 92.730 60.950 ;
        RECT 93.180 60.780 93.720 60.950 ;
        RECT 94.170 60.780 94.710 60.950 ;
        RECT 95.160 60.780 95.700 60.950 ;
        RECT 96.150 60.780 96.690 60.950 ;
        RECT 97.140 60.780 97.680 60.950 ;
        RECT 98.130 60.780 98.670 60.950 ;
        RECT 99.120 60.780 99.660 60.950 ;
        RECT 100.110 60.780 100.650 60.950 ;
        RECT 101.100 60.780 101.640 60.950 ;
        RECT 102.090 60.780 102.630 60.950 ;
        RECT 103.080 60.780 103.620 60.950 ;
        RECT 104.070 60.780 104.610 60.950 ;
        RECT 105.060 60.780 105.600 60.950 ;
        RECT 106.050 60.780 106.590 60.950 ;
        RECT 107.040 60.780 107.580 60.950 ;
        RECT 108.030 60.780 108.570 60.950 ;
        RECT 109.020 60.780 109.560 60.950 ;
        RECT 110.010 60.780 110.550 60.950 ;
        RECT 111.000 60.780 111.540 60.950 ;
        RECT 80.000 43.505 80.170 57.585 ;
        RECT 80.990 43.505 81.160 57.585 ;
        RECT 81.980 43.505 82.150 57.585 ;
        RECT 82.970 43.505 83.140 57.585 ;
        RECT 83.960 43.505 84.130 57.585 ;
        RECT 84.950 43.505 85.120 57.585 ;
        RECT 85.940 43.505 86.110 57.585 ;
        RECT 86.930 43.505 87.100 57.585 ;
        RECT 87.920 43.505 88.090 57.585 ;
        RECT 88.910 43.505 89.080 57.585 ;
        RECT 89.900 43.505 90.070 57.585 ;
        RECT 90.890 43.505 91.060 57.585 ;
        RECT 91.880 43.505 92.050 57.585 ;
        RECT 92.870 43.505 93.040 57.585 ;
        RECT 93.860 43.505 94.030 57.585 ;
        RECT 94.850 43.505 95.020 57.585 ;
        RECT 95.840 43.505 96.010 57.585 ;
        RECT 96.830 43.505 97.000 57.585 ;
        RECT 97.820 43.505 97.990 57.585 ;
        RECT 98.810 43.505 98.980 57.585 ;
        RECT 99.800 43.505 99.970 57.585 ;
        RECT 100.790 43.505 100.960 57.585 ;
        RECT 101.780 43.505 101.950 57.585 ;
        RECT 102.770 43.505 102.940 57.585 ;
        RECT 103.760 43.505 103.930 57.585 ;
        RECT 104.750 43.505 104.920 57.585 ;
        RECT 105.740 43.505 105.910 57.585 ;
        RECT 106.730 43.505 106.900 57.585 ;
        RECT 107.720 43.505 107.890 57.585 ;
        RECT 108.710 43.505 108.880 57.585 ;
        RECT 109.700 43.505 109.870 57.585 ;
        RECT 110.690 43.505 110.860 57.585 ;
        RECT 111.680 43.505 111.850 57.585 ;
        RECT 80.310 40.140 80.850 40.310 ;
        RECT 81.300 40.140 81.840 40.310 ;
        RECT 82.290 40.140 82.830 40.310 ;
        RECT 83.280 40.140 83.820 40.310 ;
        RECT 84.270 40.140 84.810 40.310 ;
        RECT 85.260 40.140 85.800 40.310 ;
        RECT 86.250 40.140 86.790 40.310 ;
        RECT 87.240 40.140 87.780 40.310 ;
        RECT 88.230 40.140 88.770 40.310 ;
        RECT 89.220 40.140 89.760 40.310 ;
        RECT 90.210 40.140 90.750 40.310 ;
        RECT 91.200 40.140 91.740 40.310 ;
        RECT 92.190 40.140 92.730 40.310 ;
        RECT 93.180 40.140 93.720 40.310 ;
        RECT 94.170 40.140 94.710 40.310 ;
        RECT 95.160 40.140 95.700 40.310 ;
        RECT 96.150 40.140 96.690 40.310 ;
        RECT 97.140 40.140 97.680 40.310 ;
        RECT 98.130 40.140 98.670 40.310 ;
        RECT 99.120 40.140 99.660 40.310 ;
        RECT 100.110 40.140 100.650 40.310 ;
        RECT 101.100 40.140 101.640 40.310 ;
        RECT 102.090 40.140 102.630 40.310 ;
        RECT 103.080 40.140 103.620 40.310 ;
        RECT 104.070 40.140 104.610 40.310 ;
        RECT 105.060 40.140 105.600 40.310 ;
        RECT 106.050 40.140 106.590 40.310 ;
        RECT 107.040 40.140 107.580 40.310 ;
        RECT 108.030 40.140 108.570 40.310 ;
        RECT 109.020 40.140 109.560 40.310 ;
        RECT 110.010 40.140 110.550 40.310 ;
        RECT 111.000 40.140 111.540 40.310 ;
        RECT 112.250 39.800 112.420 61.290 ;
        RECT 79.430 39.630 112.420 39.800 ;
      LAYER met1 ;
        RECT 1.000 220.750 8.000 222.750 ;
        RECT 7.000 196.000 8.000 220.750 ;
        RECT 3.000 194.000 74.800 196.000 ;
        RECT 6.000 191.000 72.500 193.000 ;
        RECT 16.450 189.690 61.000 189.700 ;
        RECT 13.015 189.650 61.000 189.690 ;
        RECT 12.200 189.590 61.000 189.650 ;
        RECT 12.200 189.550 62.030 189.590 ;
        RECT 64.380 189.550 65.630 189.590 ;
        RECT 67.980 189.550 69.230 189.590 ;
        RECT 69.750 189.550 70.150 189.750 ;
        RECT 12.200 189.500 16.525 189.550 ;
        RECT 12.200 187.825 12.350 189.500 ;
        RECT 13.015 189.460 16.525 189.500 ;
        RECT 19.380 189.460 20.630 189.550 ;
        RECT 60.780 189.400 70.150 189.550 ;
        RECT 13.000 189.150 13.960 189.180 ;
        RECT 14.290 189.150 15.250 189.180 ;
        RECT 15.580 189.150 16.540 189.180 ;
        RECT 17.550 189.150 17.950 189.400 ;
        RECT 60.780 189.360 62.030 189.400 ;
        RECT 64.380 189.360 65.630 189.400 ;
        RECT 67.980 189.360 69.230 189.400 ;
        RECT 19.850 189.150 20.160 189.180 ;
        RECT 13.000 189.000 32.900 189.150 ;
        RECT 61.250 189.050 61.560 189.080 ;
        RECT 64.850 189.050 65.160 189.080 ;
        RECT 68.460 189.050 68.750 189.080 ;
        RECT 13.000 188.950 13.960 189.000 ;
        RECT 14.290 188.950 15.250 189.000 ;
        RECT 15.580 188.950 16.540 189.000 ;
        RECT 19.850 188.950 20.160 189.000 ;
        RECT 32.200 188.150 32.600 188.400 ;
        RECT 14.050 188.000 19.750 188.150 ;
        RECT 12.150 180.050 12.380 187.825 ;
        RECT 14.050 187.265 14.200 188.000 ;
        RECT 16.650 187.265 16.800 188.000 ;
        RECT 12.720 180.225 12.950 187.265 ;
        RECT 14.010 180.225 14.240 187.265 ;
        RECT 15.300 180.225 15.530 187.265 ;
        RECT 16.590 180.225 16.820 187.265 ;
        RECT 12.750 180.050 12.900 180.225 ;
        RECT 15.350 180.050 15.500 180.225 ;
        RECT 12.150 179.900 15.500 180.050 ;
        RECT 12.150 179.665 12.380 179.900 ;
        RECT 17.160 179.665 17.390 187.825 ;
        RECT 19.000 179.665 19.230 187.825 ;
        RECT 19.600 187.265 19.750 188.000 ;
        RECT 20.250 188.000 32.600 188.150 ;
        RECT 20.250 187.265 20.450 188.000 ;
        RECT 19.570 180.225 19.800 187.265 ;
        RECT 20.210 187.200 20.450 187.265 ;
        RECT 20.210 180.225 20.440 187.200 ;
        RECT 20.780 179.665 21.010 187.825 ;
        RECT 32.750 182.550 32.900 189.000 ;
        RECT 60.100 188.900 65.160 189.050 ;
        RECT 33.350 188.000 33.750 188.400 ;
        RECT 60.100 184.000 60.250 188.900 ;
        RECT 61.250 188.850 61.560 188.900 ;
        RECT 64.550 187.165 64.700 188.900 ;
        RECT 64.850 188.850 65.160 188.900 ;
        RECT 68.150 188.900 68.750 189.050 ;
        RECT 68.150 187.165 68.300 188.900 ;
        RECT 68.460 188.850 68.750 188.900 ;
        RECT 68.900 187.165 69.050 189.360 ;
        RECT 69.750 189.350 70.150 189.400 ;
        RECT 58.850 183.750 59.250 184.000 ;
        RECT 59.750 183.750 60.250 184.000 ;
        RECT 58.850 183.600 60.250 183.750 ;
        RECT 42.050 183.300 59.950 183.450 ;
        RECT 33.915 182.890 37.425 183.120 ;
        RECT 40.280 182.890 41.530 183.120 ;
        RECT 42.050 182.900 42.450 183.300 ;
        RECT 44.365 182.890 47.875 183.120 ;
        RECT 50.730 182.890 51.980 183.120 ;
        RECT 33.900 182.550 34.860 182.610 ;
        RECT 35.190 182.550 36.150 182.610 ;
        RECT 36.480 182.550 37.440 182.610 ;
        RECT 40.750 182.550 41.060 182.610 ;
        RECT 44.350 182.550 45.310 182.610 ;
        RECT 45.640 182.550 46.600 182.610 ;
        RECT 46.930 182.550 47.890 182.610 ;
        RECT 51.200 182.550 51.510 182.610 ;
        RECT 32.750 182.400 51.510 182.550 ;
        RECT 33.900 182.380 34.860 182.400 ;
        RECT 35.190 182.380 36.150 182.400 ;
        RECT 36.480 182.380 37.440 182.400 ;
        RECT 37.500 181.050 37.900 181.300 ;
        RECT 34.950 180.900 37.900 181.050 ;
        RECT 34.950 180.695 35.100 180.900 ;
        RECT 37.500 180.695 37.650 180.900 ;
        RECT 12.200 178.000 12.350 179.665 ;
        RECT 13.000 178.500 13.960 178.540 ;
        RECT 14.290 178.500 15.250 178.540 ;
        RECT 15.580 178.500 16.540 178.540 ;
        RECT 17.550 178.500 17.950 178.750 ;
        RECT 19.850 178.500 20.160 178.540 ;
        RECT 13.000 178.350 20.160 178.500 ;
        RECT 13.000 178.310 13.960 178.350 ;
        RECT 14.290 178.310 15.250 178.350 ;
        RECT 15.580 178.310 16.540 178.350 ;
        RECT 19.850 178.310 20.160 178.350 ;
        RECT 13.015 178.000 16.525 178.030 ;
        RECT 19.380 178.000 20.630 178.030 ;
        RECT 20.800 178.000 20.950 179.665 ;
        RECT 33.050 178.000 33.280 179.580 ;
        RECT 12.200 177.850 33.280 178.000 ;
        RECT 12.200 169.335 12.350 177.850 ;
        RECT 13.015 177.800 16.525 177.850 ;
        RECT 19.380 177.800 20.630 177.850 ;
        RECT 21.150 176.550 31.750 176.700 ;
        RECT 13.015 176.000 16.525 176.230 ;
        RECT 19.380 176.000 20.630 176.230 ;
        RECT 13.000 175.700 13.960 175.720 ;
        RECT 14.290 175.700 15.250 175.720 ;
        RECT 15.580 175.700 16.540 175.720 ;
        RECT 17.550 175.700 17.950 175.950 ;
        RECT 19.850 175.700 20.160 175.720 ;
        RECT 13.000 175.550 21.000 175.700 ;
        RECT 13.000 175.490 13.960 175.550 ;
        RECT 14.290 175.490 15.250 175.550 ;
        RECT 15.580 175.490 16.540 175.550 ;
        RECT 16.600 174.150 17.000 174.400 ;
        RECT 14.050 174.000 17.000 174.150 ;
        RECT 14.050 173.805 14.200 174.000 ;
        RECT 16.650 173.805 16.800 174.000 ;
        RECT 12.150 166.550 12.380 169.335 ;
        RECT 12.720 166.765 12.950 173.805 ;
        RECT 14.010 166.765 14.240 173.805 ;
        RECT 15.300 166.765 15.530 173.805 ;
        RECT 16.590 166.765 16.820 173.805 ;
        RECT 12.750 166.550 12.900 166.765 ;
        RECT 15.350 166.550 15.500 166.765 ;
        RECT 12.150 166.400 15.500 166.550 ;
        RECT 12.150 155.350 12.380 166.400 ;
        RECT 13.000 165.050 13.960 165.080 ;
        RECT 14.290 165.050 15.250 165.080 ;
        RECT 15.580 165.050 16.540 165.080 ;
        RECT 13.000 164.900 16.600 165.050 ;
        RECT 13.000 164.850 17.000 164.900 ;
        RECT 13.050 164.540 17.000 164.850 ;
        RECT 13.000 164.500 17.000 164.540 ;
        RECT 13.000 164.350 16.600 164.500 ;
        RECT 13.000 164.310 13.960 164.350 ;
        RECT 14.290 164.310 15.250 164.350 ;
        RECT 15.580 164.310 16.540 164.350 ;
        RECT 16.600 162.950 17.000 163.200 ;
        RECT 14.050 162.800 17.000 162.950 ;
        RECT 14.050 162.625 14.200 162.800 ;
        RECT 16.650 162.625 16.800 162.800 ;
        RECT 12.720 155.585 12.950 162.625 ;
        RECT 14.010 155.585 14.240 162.625 ;
        RECT 15.300 155.585 15.530 162.625 ;
        RECT 16.590 155.585 16.820 162.625 ;
        RECT 12.750 155.350 12.900 155.585 ;
        RECT 15.350 155.350 15.500 155.585 ;
        RECT 12.150 155.200 15.500 155.350 ;
        RECT 12.150 144.200 12.380 155.200 ;
        RECT 13.000 153.850 13.960 153.900 ;
        RECT 14.290 153.850 15.250 153.900 ;
        RECT 15.580 153.850 16.540 153.900 ;
        RECT 13.000 153.750 16.600 153.850 ;
        RECT 13.000 153.670 17.000 153.750 ;
        RECT 13.050 153.360 17.000 153.670 ;
        RECT 13.000 153.350 17.000 153.360 ;
        RECT 13.000 153.200 16.600 153.350 ;
        RECT 13.000 153.130 13.960 153.200 ;
        RECT 14.290 153.130 15.250 153.200 ;
        RECT 15.580 153.130 16.540 153.200 ;
        RECT 16.600 151.850 17.000 152.100 ;
        RECT 14.050 151.700 17.000 151.850 ;
        RECT 14.050 151.445 14.200 151.700 ;
        RECT 16.650 151.445 16.800 151.700 ;
        RECT 12.720 144.405 12.950 151.445 ;
        RECT 14.010 144.405 14.240 151.445 ;
        RECT 15.300 144.405 15.530 151.445 ;
        RECT 16.590 144.405 16.820 151.445 ;
        RECT 12.750 144.200 12.900 144.405 ;
        RECT 15.350 144.200 15.500 144.405 ;
        RECT 12.150 144.050 15.500 144.200 ;
        RECT 12.150 137.695 12.380 144.050 ;
        RECT 13.000 142.700 13.960 142.720 ;
        RECT 14.290 142.700 15.250 142.720 ;
        RECT 15.580 142.700 16.540 142.720 ;
        RECT 13.000 142.550 16.600 142.700 ;
        RECT 13.000 142.490 17.000 142.550 ;
        RECT 13.050 142.180 17.000 142.490 ;
        RECT 13.000 142.150 17.000 142.180 ;
        RECT 13.000 142.000 16.600 142.150 ;
        RECT 13.000 141.950 13.960 142.000 ;
        RECT 14.290 141.950 15.250 142.000 ;
        RECT 15.580 141.950 16.540 142.000 ;
        RECT 16.600 140.600 17.000 140.850 ;
        RECT 14.050 140.450 17.000 140.600 ;
        RECT 14.050 140.265 14.200 140.450 ;
        RECT 16.650 140.265 16.800 140.450 ;
        RECT 12.200 133.000 12.350 137.695 ;
        RECT 12.720 133.225 12.950 140.265 ;
        RECT 14.010 133.225 14.240 140.265 ;
        RECT 15.300 133.225 15.530 140.265 ;
        RECT 16.590 133.225 16.820 140.265 ;
        RECT 17.160 137.695 17.390 169.335 ;
        RECT 17.550 165.050 17.700 175.550 ;
        RECT 19.850 175.490 20.160 175.550 ;
        RECT 20.600 175.300 21.000 175.550 ;
        RECT 17.850 173.850 18.250 174.250 ;
        RECT 19.400 174.000 19.800 174.400 ;
        RECT 17.550 164.650 17.950 165.050 ;
        RECT 17.550 153.900 17.700 164.650 ;
        RECT 18.100 163.350 18.250 173.850 ;
        RECT 19.600 173.805 19.750 174.000 ;
        RECT 18.100 162.950 18.500 163.350 ;
        RECT 17.550 153.500 17.950 153.900 ;
        RECT 17.550 142.700 17.700 153.500 ;
        RECT 18.100 152.250 18.250 162.950 ;
        RECT 18.100 151.850 18.500 152.250 ;
        RECT 17.550 142.300 17.950 142.700 ;
        RECT 12.750 133.000 12.900 133.225 ;
        RECT 15.350 133.000 15.500 133.225 ;
        RECT 12.200 132.850 15.500 133.000 ;
        RECT 12.200 131.000 12.350 132.850 ;
        RECT 17.550 131.900 17.700 142.300 ;
        RECT 18.100 141.000 18.250 151.850 ;
        RECT 18.100 140.600 18.500 141.000 ;
        RECT 19.000 137.695 19.230 169.335 ;
        RECT 19.570 166.765 19.800 173.805 ;
        RECT 20.210 173.750 20.440 173.805 ;
        RECT 21.150 173.750 21.300 176.550 ;
        RECT 23.465 176.150 26.975 176.380 ;
        RECT 29.830 176.150 31.080 176.380 ;
        RECT 23.450 175.850 24.410 175.870 ;
        RECT 24.740 175.850 25.700 175.870 ;
        RECT 26.030 175.850 26.990 175.870 ;
        RECT 30.300 175.850 30.610 175.870 ;
        RECT 22.050 175.700 30.610 175.850 ;
        RECT 22.050 175.450 22.450 175.700 ;
        RECT 23.450 175.640 24.410 175.700 ;
        RECT 24.740 175.640 25.700 175.700 ;
        RECT 26.030 175.640 26.990 175.700 ;
        RECT 27.050 174.300 27.450 174.550 ;
        RECT 24.500 174.150 27.450 174.300 ;
        RECT 24.500 173.955 24.650 174.150 ;
        RECT 27.100 173.955 27.250 174.150 ;
        RECT 20.210 173.600 21.300 173.750 ;
        RECT 20.210 167.000 20.440 173.600 ;
        RECT 20.210 166.765 20.500 167.000 ;
        RECT 19.850 165.050 20.160 165.080 ;
        RECT 19.800 164.900 20.160 165.050 ;
        RECT 19.400 164.850 20.160 164.900 ;
        RECT 19.400 164.540 20.100 164.850 ;
        RECT 19.400 164.500 20.160 164.540 ;
        RECT 19.800 164.350 20.160 164.500 ;
        RECT 19.850 164.310 20.160 164.350 ;
        RECT 19.400 162.800 19.800 163.200 ;
        RECT 19.600 162.625 19.750 162.800 ;
        RECT 20.350 162.625 20.500 166.765 ;
        RECT 19.570 155.585 19.800 162.625 ;
        RECT 20.210 162.400 20.500 162.625 ;
        RECT 20.210 155.800 20.440 162.400 ;
        RECT 20.210 155.585 20.500 155.800 ;
        RECT 19.850 153.850 20.160 153.900 ;
        RECT 19.800 153.750 20.160 153.850 ;
        RECT 19.400 153.670 20.160 153.750 ;
        RECT 19.400 153.360 20.100 153.670 ;
        RECT 19.400 153.350 20.160 153.360 ;
        RECT 19.800 153.150 20.160 153.350 ;
        RECT 19.850 153.130 20.160 153.150 ;
        RECT 19.400 151.700 19.800 152.100 ;
        RECT 19.600 151.445 19.750 151.700 ;
        RECT 20.350 151.445 20.500 155.585 ;
        RECT 19.570 144.405 19.800 151.445 ;
        RECT 20.210 151.200 20.500 151.445 ;
        RECT 20.210 144.600 20.440 151.200 ;
        RECT 20.210 144.405 20.500 144.600 ;
        RECT 19.850 142.700 20.160 142.720 ;
        RECT 19.800 142.550 20.160 142.700 ;
        RECT 19.400 142.490 20.160 142.550 ;
        RECT 19.400 142.180 20.100 142.490 ;
        RECT 19.400 142.150 20.160 142.180 ;
        RECT 19.800 142.000 20.160 142.150 ;
        RECT 19.850 141.950 20.160 142.000 ;
        RECT 19.400 140.450 19.800 140.850 ;
        RECT 19.600 140.265 19.750 140.450 ;
        RECT 20.350 140.265 20.500 144.405 ;
        RECT 19.570 133.225 19.800 140.265 ;
        RECT 20.210 140.050 20.500 140.265 ;
        RECT 20.210 133.225 20.440 140.050 ;
        RECT 20.780 137.695 21.010 169.335 ;
        RECT 22.600 166.750 22.830 169.485 ;
        RECT 23.170 166.915 23.400 173.955 ;
        RECT 24.460 166.915 24.690 173.955 ;
        RECT 25.750 166.915 25.980 173.955 ;
        RECT 27.040 166.915 27.270 173.955 ;
        RECT 23.200 166.750 23.350 166.915 ;
        RECT 25.800 166.750 25.950 166.915 ;
        RECT 22.600 166.600 25.950 166.750 ;
        RECT 22.600 155.550 22.830 166.600 ;
        RECT 23.450 165.200 24.410 165.230 ;
        RECT 24.740 165.200 25.700 165.230 ;
        RECT 26.030 165.200 26.990 165.230 ;
        RECT 23.450 165.050 27.050 165.200 ;
        RECT 23.450 165.000 27.450 165.050 ;
        RECT 23.500 164.690 27.450 165.000 ;
        RECT 23.450 164.650 27.450 164.690 ;
        RECT 23.450 164.500 27.050 164.650 ;
        RECT 23.450 164.460 24.410 164.500 ;
        RECT 24.740 164.460 25.700 164.500 ;
        RECT 26.030 164.460 26.990 164.500 ;
        RECT 27.050 163.100 27.450 163.350 ;
        RECT 24.500 162.950 27.450 163.100 ;
        RECT 24.500 162.775 24.650 162.950 ;
        RECT 27.050 162.775 27.200 162.950 ;
        RECT 23.170 155.735 23.400 162.775 ;
        RECT 24.460 155.735 24.690 162.775 ;
        RECT 25.750 155.735 25.980 162.775 ;
        RECT 27.040 155.735 27.270 162.775 ;
        RECT 23.200 155.550 23.350 155.735 ;
        RECT 25.800 155.550 25.950 155.735 ;
        RECT 22.600 155.400 25.950 155.550 ;
        RECT 22.600 144.400 22.830 155.400 ;
        RECT 23.450 154.000 24.410 154.050 ;
        RECT 24.740 154.000 25.700 154.050 ;
        RECT 26.030 154.000 26.990 154.050 ;
        RECT 23.450 153.850 27.050 154.000 ;
        RECT 23.450 153.820 27.450 153.850 ;
        RECT 23.500 153.510 27.450 153.820 ;
        RECT 23.450 153.450 27.450 153.510 ;
        RECT 23.450 153.300 27.050 153.450 ;
        RECT 23.450 153.280 24.410 153.300 ;
        RECT 24.740 153.280 25.700 153.300 ;
        RECT 26.030 153.280 26.990 153.300 ;
        RECT 27.050 151.950 27.450 152.200 ;
        RECT 24.500 151.800 27.450 151.950 ;
        RECT 24.500 151.595 24.650 151.800 ;
        RECT 27.050 151.595 27.200 151.800 ;
        RECT 23.170 144.555 23.400 151.595 ;
        RECT 24.460 144.555 24.690 151.595 ;
        RECT 25.750 144.555 25.980 151.595 ;
        RECT 27.040 144.555 27.270 151.595 ;
        RECT 23.200 144.400 23.350 144.555 ;
        RECT 25.800 144.400 25.950 144.555 ;
        RECT 22.600 144.250 25.950 144.400 ;
        RECT 22.600 137.845 22.830 144.250 ;
        RECT 23.450 142.850 24.410 142.870 ;
        RECT 24.740 142.850 25.700 142.870 ;
        RECT 26.030 142.850 26.990 142.870 ;
        RECT 23.450 142.650 27.050 142.850 ;
        RECT 23.450 142.640 27.450 142.650 ;
        RECT 23.550 142.330 27.450 142.640 ;
        RECT 23.450 142.250 27.450 142.330 ;
        RECT 23.450 142.150 27.050 142.250 ;
        RECT 23.450 142.100 24.410 142.150 ;
        RECT 24.740 142.100 25.700 142.150 ;
        RECT 26.030 142.100 26.990 142.150 ;
        RECT 27.050 140.750 27.450 141.000 ;
        RECT 24.500 140.600 27.450 140.750 ;
        RECT 24.500 140.415 24.650 140.600 ;
        RECT 27.050 140.415 27.200 140.600 ;
        RECT 13.000 131.500 13.960 131.540 ;
        RECT 14.290 131.500 15.250 131.540 ;
        RECT 15.580 131.500 16.540 131.540 ;
        RECT 17.550 131.500 17.950 131.900 ;
        RECT 19.850 131.500 20.160 131.540 ;
        RECT 13.000 131.350 20.160 131.500 ;
        RECT 13.000 131.310 13.960 131.350 ;
        RECT 14.290 131.310 15.250 131.350 ;
        RECT 15.580 131.310 16.540 131.350 ;
        RECT 19.850 131.310 20.160 131.350 ;
        RECT 20.800 131.150 20.950 137.695 ;
        RECT 22.650 133.200 22.800 137.845 ;
        RECT 23.170 133.375 23.400 140.415 ;
        RECT 24.460 133.375 24.690 140.415 ;
        RECT 25.750 133.375 25.980 140.415 ;
        RECT 27.040 133.375 27.270 140.415 ;
        RECT 27.610 137.845 27.840 169.485 ;
        RECT 28.000 165.200 28.150 175.700 ;
        RECT 30.300 175.640 30.610 175.700 ;
        RECT 28.900 174.300 29.300 174.700 ;
        RECT 28.000 164.800 28.400 165.200 ;
        RECT 28.000 154.000 28.150 164.800 ;
        RECT 29.150 163.500 29.300 174.300 ;
        RECT 29.850 174.150 30.250 174.550 ;
        RECT 30.100 173.955 30.250 174.150 ;
        RECT 28.900 163.100 29.300 163.500 ;
        RECT 28.000 153.600 28.400 154.000 ;
        RECT 28.000 142.800 28.150 153.600 ;
        RECT 29.150 152.350 29.300 163.100 ;
        RECT 28.900 151.950 29.300 152.350 ;
        RECT 28.000 142.400 28.400 142.800 ;
        RECT 23.200 133.200 23.350 133.375 ;
        RECT 25.800 133.200 25.950 133.375 ;
        RECT 22.650 133.050 25.950 133.200 ;
        RECT 22.650 131.150 22.800 133.050 ;
        RECT 23.450 131.650 24.410 131.690 ;
        RECT 24.740 131.650 25.700 131.690 ;
        RECT 26.030 131.650 26.990 131.690 ;
        RECT 28.000 131.650 28.150 142.400 ;
        RECT 29.150 141.150 29.300 151.950 ;
        RECT 28.900 140.750 29.300 141.150 ;
        RECT 29.450 137.845 29.680 169.485 ;
        RECT 30.020 166.915 30.250 173.955 ;
        RECT 30.660 169.800 30.890 173.955 ;
        RECT 31.050 169.800 31.450 170.050 ;
        RECT 30.660 169.650 31.450 169.800 ;
        RECT 30.660 167.100 30.890 169.650 ;
        RECT 30.660 166.915 30.950 167.100 ;
        RECT 30.300 165.200 30.610 165.230 ;
        RECT 30.250 165.050 30.610 165.200 ;
        RECT 29.850 165.000 30.610 165.050 ;
        RECT 29.850 164.690 30.600 165.000 ;
        RECT 29.850 164.650 30.610 164.690 ;
        RECT 30.250 164.500 30.610 164.650 ;
        RECT 30.300 164.460 30.610 164.500 ;
        RECT 29.850 162.950 30.250 163.350 ;
        RECT 30.100 162.775 30.250 162.950 ;
        RECT 30.800 162.775 30.950 166.915 ;
        RECT 30.020 155.735 30.250 162.775 ;
        RECT 30.660 162.550 30.950 162.775 ;
        RECT 30.660 155.950 30.890 162.550 ;
        RECT 30.660 155.735 30.950 155.950 ;
        RECT 30.300 154.000 30.610 154.050 ;
        RECT 30.250 153.850 30.610 154.000 ;
        RECT 29.850 153.820 30.610 153.850 ;
        RECT 29.850 153.510 30.550 153.820 ;
        RECT 29.850 153.450 30.610 153.510 ;
        RECT 30.250 153.300 30.610 153.450 ;
        RECT 30.300 153.280 30.610 153.300 ;
        RECT 29.850 151.800 30.250 152.200 ;
        RECT 30.100 151.595 30.250 151.800 ;
        RECT 30.800 151.595 30.950 155.735 ;
        RECT 30.020 144.555 30.250 151.595 ;
        RECT 30.660 151.400 30.950 151.595 ;
        RECT 30.660 144.750 30.890 151.400 ;
        RECT 30.660 144.555 30.950 144.750 ;
        RECT 30.300 142.850 30.610 142.870 ;
        RECT 30.250 142.650 30.610 142.850 ;
        RECT 29.850 142.640 30.610 142.650 ;
        RECT 29.850 142.330 30.550 142.640 ;
        RECT 29.850 142.250 30.610 142.330 ;
        RECT 30.250 142.100 30.610 142.250 ;
        RECT 29.850 140.600 30.250 141.000 ;
        RECT 30.100 140.415 30.250 140.600 ;
        RECT 30.800 140.415 30.950 144.555 ;
        RECT 30.020 133.375 30.250 140.415 ;
        RECT 30.660 140.200 30.950 140.415 ;
        RECT 30.660 133.375 30.890 140.200 ;
        RECT 31.230 137.845 31.460 169.485 ;
        RECT 31.600 159.300 31.750 176.550 ;
        RECT 33.050 173.450 33.280 177.850 ;
        RECT 33.620 173.655 33.850 180.695 ;
        RECT 34.910 173.655 35.140 180.695 ;
        RECT 36.200 173.655 36.430 180.695 ;
        RECT 37.490 173.655 37.720 180.695 ;
        RECT 33.650 173.450 33.800 173.655 ;
        RECT 36.250 173.450 36.400 173.655 ;
        RECT 33.050 173.300 36.400 173.450 ;
        RECT 33.050 163.590 33.280 173.300 ;
        RECT 33.900 171.950 34.860 171.970 ;
        RECT 35.190 171.950 36.150 171.970 ;
        RECT 36.480 171.950 37.440 171.970 ;
        RECT 33.900 171.800 37.500 171.950 ;
        RECT 33.900 171.740 37.900 171.800 ;
        RECT 33.950 171.430 37.900 171.740 ;
        RECT 33.900 171.400 37.900 171.430 ;
        RECT 33.900 171.250 37.500 171.400 ;
        RECT 33.900 171.200 34.860 171.250 ;
        RECT 35.190 171.200 36.150 171.250 ;
        RECT 36.480 171.200 37.440 171.250 ;
        RECT 37.500 169.850 37.900 170.100 ;
        RECT 34.950 169.700 37.900 169.850 ;
        RECT 34.950 169.515 35.100 169.700 ;
        RECT 37.500 169.515 37.650 169.700 ;
        RECT 33.050 162.300 33.200 163.590 ;
        RECT 33.620 162.475 33.850 169.515 ;
        RECT 34.910 162.475 35.140 169.515 ;
        RECT 36.200 162.475 36.430 169.515 ;
        RECT 37.490 162.475 37.720 169.515 ;
        RECT 38.060 163.590 38.290 179.580 ;
        RECT 38.450 171.950 38.600 182.400 ;
        RECT 40.750 182.380 41.060 182.400 ;
        RECT 44.350 182.380 45.310 182.400 ;
        RECT 45.640 182.380 46.600 182.400 ;
        RECT 46.930 182.380 47.890 182.400 ;
        RECT 39.350 181.050 39.750 181.450 ;
        RECT 38.450 171.550 38.850 171.950 ;
        RECT 33.650 162.300 33.800 162.475 ;
        RECT 36.250 162.300 36.400 162.475 ;
        RECT 33.050 162.150 36.400 162.300 ;
        RECT 33.050 160.250 33.200 162.150 ;
        RECT 33.900 160.750 34.860 160.790 ;
        RECT 35.190 160.750 36.150 160.790 ;
        RECT 36.480 160.750 37.440 160.790 ;
        RECT 38.450 160.750 38.600 171.550 ;
        RECT 39.600 170.250 39.750 181.050 ;
        RECT 40.300 180.900 40.700 181.300 ;
        RECT 47.950 181.050 48.350 181.300 ;
        RECT 45.400 180.900 48.350 181.050 ;
        RECT 40.500 180.695 40.650 180.900 ;
        RECT 39.350 169.850 39.750 170.250 ;
        RECT 39.900 163.590 40.130 179.580 ;
        RECT 40.470 173.655 40.700 180.695 ;
        RECT 41.110 180.650 41.340 180.695 ;
        RECT 42.050 180.650 42.450 180.900 ;
        RECT 45.400 180.695 45.550 180.900 ;
        RECT 47.950 180.695 48.100 180.900 ;
        RECT 41.110 180.500 42.450 180.650 ;
        RECT 41.110 173.850 41.340 180.500 ;
        RECT 41.110 173.655 41.400 173.850 ;
        RECT 40.750 171.950 41.060 171.970 ;
        RECT 40.700 171.800 41.060 171.950 ;
        RECT 40.300 171.740 41.060 171.800 ;
        RECT 40.300 171.430 41.000 171.740 ;
        RECT 40.300 171.400 41.060 171.430 ;
        RECT 40.700 171.250 41.060 171.400 ;
        RECT 40.750 171.200 41.060 171.250 ;
        RECT 40.300 169.700 40.700 170.100 ;
        RECT 40.500 169.515 40.650 169.700 ;
        RECT 41.250 169.515 41.400 173.655 ;
        RECT 40.470 162.475 40.700 169.515 ;
        RECT 41.110 169.300 41.400 169.515 ;
        RECT 41.110 162.475 41.340 169.300 ;
        RECT 41.680 163.590 41.910 179.580 ;
        RECT 43.500 173.450 43.730 179.580 ;
        RECT 44.070 173.655 44.300 180.695 ;
        RECT 45.360 173.655 45.590 180.695 ;
        RECT 46.650 173.655 46.880 180.695 ;
        RECT 47.940 173.655 48.170 180.695 ;
        RECT 44.100 173.450 44.250 173.655 ;
        RECT 46.700 173.450 46.850 173.655 ;
        RECT 43.500 173.300 46.850 173.450 ;
        RECT 43.500 163.590 43.730 173.300 ;
        RECT 44.350 171.950 45.310 171.970 ;
        RECT 45.640 171.950 46.600 171.970 ;
        RECT 46.930 171.950 47.890 171.970 ;
        RECT 44.350 171.800 47.950 171.950 ;
        RECT 44.350 171.740 48.350 171.800 ;
        RECT 44.400 171.430 48.350 171.740 ;
        RECT 44.350 171.400 48.350 171.430 ;
        RECT 44.350 171.250 47.950 171.400 ;
        RECT 44.350 171.200 45.310 171.250 ;
        RECT 45.640 171.200 46.600 171.250 ;
        RECT 46.930 171.200 47.890 171.250 ;
        RECT 47.950 169.850 48.350 170.100 ;
        RECT 45.400 169.700 48.350 169.850 ;
        RECT 45.400 169.515 45.550 169.700 ;
        RECT 48.000 169.515 48.150 169.700 ;
        RECT 40.750 160.750 41.060 160.790 ;
        RECT 33.900 160.600 41.060 160.750 ;
        RECT 33.900 160.560 34.860 160.600 ;
        RECT 35.190 160.560 36.150 160.600 ;
        RECT 36.480 160.560 37.440 160.600 ;
        RECT 40.750 160.560 41.060 160.600 ;
        RECT 33.915 160.250 37.425 160.280 ;
        RECT 40.280 160.250 41.530 160.280 ;
        RECT 41.750 160.250 41.900 163.590 ;
        RECT 43.550 162.300 43.700 163.590 ;
        RECT 44.070 162.475 44.300 169.515 ;
        RECT 45.360 162.475 45.590 169.515 ;
        RECT 46.650 162.475 46.880 169.515 ;
        RECT 47.940 162.475 48.170 169.515 ;
        RECT 48.510 163.590 48.740 179.580 ;
        RECT 48.900 171.950 49.050 182.400 ;
        RECT 51.200 182.380 51.510 182.400 ;
        RECT 49.800 181.050 50.200 181.450 ;
        RECT 48.900 171.550 49.450 171.950 ;
        RECT 44.100 162.300 44.250 162.475 ;
        RECT 46.700 162.300 46.850 162.475 ;
        RECT 43.550 162.150 46.850 162.300 ;
        RECT 43.550 160.250 43.700 162.150 ;
        RECT 44.350 160.750 45.310 160.790 ;
        RECT 45.640 160.750 46.600 160.790 ;
        RECT 46.930 160.750 47.890 160.790 ;
        RECT 48.900 160.750 49.050 171.550 ;
        RECT 50.050 170.250 50.200 181.050 ;
        RECT 50.750 180.900 51.150 181.300 ;
        RECT 50.950 180.695 51.100 180.900 ;
        RECT 49.800 169.850 50.200 170.250 ;
        RECT 50.350 163.590 50.580 179.580 ;
        RECT 50.920 173.655 51.150 180.695 ;
        RECT 51.560 180.650 51.790 180.695 ;
        RECT 51.560 180.500 52.650 180.650 ;
        RECT 51.560 173.850 51.790 180.500 ;
        RECT 51.560 173.655 51.850 173.850 ;
        RECT 51.200 171.950 51.510 171.970 ;
        RECT 51.150 171.800 51.510 171.950 ;
        RECT 50.750 171.740 51.510 171.800 ;
        RECT 50.750 171.430 51.450 171.740 ;
        RECT 50.750 171.400 51.510 171.430 ;
        RECT 51.150 171.250 51.510 171.400 ;
        RECT 51.200 171.200 51.510 171.250 ;
        RECT 50.750 169.700 51.150 170.100 ;
        RECT 50.950 169.515 51.100 169.700 ;
        RECT 51.700 169.515 51.850 173.655 ;
        RECT 50.920 162.475 51.150 169.515 ;
        RECT 51.560 169.300 51.850 169.515 ;
        RECT 51.560 162.475 51.790 169.300 ;
        RECT 52.130 163.590 52.360 179.580 ;
        RECT 51.200 160.750 51.510 160.790 ;
        RECT 44.350 160.600 51.510 160.750 ;
        RECT 44.350 160.560 45.310 160.600 ;
        RECT 45.640 160.560 46.600 160.600 ;
        RECT 46.930 160.560 47.890 160.600 ;
        RECT 51.200 160.560 51.510 160.600 ;
        RECT 48.900 160.300 50.200 160.450 ;
        RECT 44.365 160.250 47.875 160.280 ;
        RECT 48.900 160.250 49.050 160.300 ;
        RECT 33.050 160.100 49.050 160.250 ;
        RECT 50.050 160.250 50.200 160.300 ;
        RECT 50.730 160.250 51.980 160.280 ;
        RECT 52.200 160.250 52.350 163.590 ;
        RECT 33.915 160.050 37.425 160.100 ;
        RECT 40.280 160.050 41.530 160.100 ;
        RECT 44.365 160.050 47.875 160.100 ;
        RECT 49.200 159.900 49.600 160.150 ;
        RECT 50.050 160.100 52.350 160.250 ;
        RECT 50.730 160.050 51.980 160.100 ;
        RECT 34.500 159.750 49.600 159.900 ;
        RECT 52.200 159.750 52.350 160.100 ;
        RECT 52.500 160.050 52.650 180.500 ;
        RECT 59.800 177.550 59.950 183.300 ;
        RECT 60.100 178.400 60.250 183.600 ;
        RECT 60.970 180.350 61.200 187.165 ;
        RECT 60.650 180.200 61.200 180.350 ;
        RECT 60.650 179.050 60.800 180.200 ;
        RECT 60.970 180.125 61.200 180.200 ;
        RECT 61.610 180.350 61.840 187.165 ;
        RECT 64.550 186.950 64.800 187.165 ;
        RECT 64.570 180.350 64.800 186.950 ;
        RECT 61.610 180.200 62.700 180.350 ;
        RECT 61.610 180.125 61.840 180.200 ;
        RECT 60.400 178.650 60.800 179.050 ;
        RECT 61.250 178.400 61.560 178.440 ;
        RECT 60.100 178.250 61.560 178.400 ;
        RECT 61.250 178.210 61.560 178.250 ;
        RECT 62.550 177.950 62.700 180.200 ;
        RECT 64.550 180.125 64.800 180.350 ;
        RECT 65.210 187.100 65.440 187.165 ;
        RECT 68.150 187.100 68.400 187.165 ;
        RECT 65.210 186.950 68.400 187.100 ;
        RECT 65.210 180.125 65.440 186.950 ;
        RECT 68.170 180.350 68.400 186.950 ;
        RECT 68.150 180.125 68.400 180.350 ;
        RECT 68.810 186.950 69.050 187.165 ;
        RECT 68.810 180.125 69.040 186.950 ;
        RECT 64.550 178.400 64.700 180.125 ;
        RECT 64.850 178.400 65.160 178.440 ;
        RECT 64.550 178.250 65.160 178.400 ;
        RECT 68.150 178.400 68.300 180.125 ;
        RECT 68.460 178.400 68.750 178.440 ;
        RECT 68.150 178.250 68.750 178.400 ;
        RECT 64.850 178.210 65.160 178.250 ;
        RECT 68.460 178.210 68.750 178.250 ;
        RECT 62.550 177.550 62.950 177.950 ;
        RECT 59.800 177.400 62.700 177.550 ;
        RECT 59.800 166.150 59.950 177.400 ;
        RECT 59.800 166.000 60.750 166.150 ;
        RECT 60.350 165.750 60.750 166.000 ;
        RECT 67.980 165.600 69.230 165.650 ;
        RECT 70.500 165.600 72.500 191.000 ;
        RECT 72.800 188.300 74.800 194.000 ;
        RECT 75.450 189.050 75.760 189.060 ;
        RECT 76.090 189.050 76.400 189.060 ;
        RECT 76.730 189.050 77.040 189.060 ;
        RECT 77.370 189.050 77.680 189.060 ;
        RECT 78.010 189.050 78.320 189.060 ;
        RECT 78.650 189.050 78.960 189.060 ;
        RECT 79.290 189.050 79.600 189.060 ;
        RECT 79.930 189.050 80.240 189.060 ;
        RECT 80.570 189.050 80.880 189.060 ;
        RECT 81.210 189.050 81.520 189.060 ;
        RECT 81.850 189.050 82.160 189.060 ;
        RECT 75.450 188.850 82.950 189.050 ;
        RECT 75.450 188.830 75.760 188.850 ;
        RECT 76.090 188.830 76.400 188.850 ;
        RECT 76.730 188.830 77.040 188.850 ;
        RECT 77.370 188.830 77.680 188.850 ;
        RECT 78.010 188.830 78.320 188.850 ;
        RECT 78.650 188.830 78.960 188.850 ;
        RECT 79.290 188.830 79.600 188.850 ;
        RECT 79.930 188.830 80.240 188.850 ;
        RECT 80.570 188.830 80.880 188.850 ;
        RECT 81.210 188.830 81.520 188.850 ;
        RECT 81.850 188.830 82.160 188.850 ;
        RECT 82.550 188.650 82.950 188.850 ;
        RECT 72.800 187.300 81.800 188.300 ;
        RECT 72.800 186.030 74.800 187.300 ;
        RECT 75.200 187.145 75.400 187.300 ;
        RECT 76.450 187.145 76.650 187.300 ;
        RECT 77.750 187.145 77.950 187.300 ;
        RECT 79.000 187.145 79.200 187.300 ;
        RECT 80.300 187.145 80.500 187.300 ;
        RECT 81.600 187.145 81.800 187.300 ;
        RECT 72.800 170.040 74.830 186.030 ;
        RECT 75.170 180.105 75.400 187.145 ;
        RECT 75.810 180.150 76.040 187.145 ;
        RECT 75.800 180.105 76.040 180.150 ;
        RECT 76.450 180.105 76.680 187.145 ;
        RECT 77.090 180.105 77.320 187.145 ;
        RECT 77.730 180.105 77.960 187.145 ;
        RECT 78.370 180.105 78.600 187.145 ;
        RECT 79.000 187.100 79.240 187.145 ;
        RECT 79.010 180.105 79.240 187.100 ;
        RECT 79.650 180.105 79.880 187.145 ;
        RECT 80.290 180.105 80.520 187.145 ;
        RECT 80.930 180.105 81.160 187.145 ;
        RECT 81.570 180.105 81.800 187.145 ;
        RECT 82.210 180.150 82.440 187.145 ;
        RECT 82.200 180.105 82.440 180.150 ;
        RECT 75.800 179.950 76.000 180.105 ;
        RECT 77.100 179.950 77.300 180.105 ;
        RECT 78.400 179.950 78.600 180.105 ;
        RECT 79.650 179.950 79.850 180.105 ;
        RECT 80.950 179.950 81.150 180.105 ;
        RECT 82.200 179.950 82.400 180.105 ;
        RECT 75.800 178.950 87.100 179.950 ;
        RECT 75.450 178.400 75.760 178.420 ;
        RECT 76.090 178.400 76.400 178.420 ;
        RECT 76.730 178.400 77.040 178.420 ;
        RECT 77.370 178.400 77.680 178.420 ;
        RECT 78.010 178.400 78.320 178.420 ;
        RECT 78.650 178.400 78.960 178.420 ;
        RECT 79.290 178.400 79.600 178.420 ;
        RECT 79.930 178.400 80.240 178.420 ;
        RECT 80.570 178.400 80.880 178.420 ;
        RECT 81.210 178.400 81.520 178.420 ;
        RECT 81.850 178.400 82.160 178.420 ;
        RECT 75.450 178.250 82.550 178.400 ;
        RECT 75.450 178.190 82.950 178.250 ;
        RECT 75.500 177.880 82.950 178.190 ;
        RECT 75.450 177.850 82.950 177.880 ;
        RECT 75.450 177.700 82.550 177.850 ;
        RECT 75.450 177.650 75.760 177.700 ;
        RECT 76.090 177.650 76.400 177.700 ;
        RECT 76.730 177.650 77.040 177.700 ;
        RECT 77.370 177.650 77.680 177.700 ;
        RECT 78.010 177.650 78.320 177.700 ;
        RECT 78.650 177.650 78.960 177.700 ;
        RECT 79.290 177.650 79.600 177.700 ;
        RECT 79.930 177.650 80.240 177.700 ;
        RECT 80.570 177.650 80.880 177.700 ;
        RECT 81.210 177.650 81.520 177.700 ;
        RECT 81.850 177.650 82.160 177.700 ;
        RECT 85.100 177.150 87.100 178.950 ;
        RECT 75.800 176.150 87.100 177.150 ;
        RECT 75.800 175.965 76.000 176.150 ;
        RECT 77.100 175.965 77.300 176.150 ;
        RECT 78.350 175.965 78.550 176.150 ;
        RECT 79.650 175.965 79.850 176.150 ;
        RECT 80.950 175.965 81.150 176.150 ;
        RECT 82.200 175.965 82.400 176.150 ;
        RECT 72.800 168.750 74.800 170.040 ;
        RECT 75.170 168.925 75.400 175.965 ;
        RECT 75.800 175.900 76.040 175.965 ;
        RECT 75.810 168.925 76.040 175.900 ;
        RECT 76.450 168.925 76.680 175.965 ;
        RECT 77.090 168.925 77.320 175.965 ;
        RECT 77.730 168.925 77.960 175.965 ;
        RECT 78.350 175.900 78.600 175.965 ;
        RECT 78.370 168.925 78.600 175.900 ;
        RECT 79.010 169.000 79.240 175.965 ;
        RECT 79.000 168.925 79.240 169.000 ;
        RECT 79.650 168.925 79.880 175.965 ;
        RECT 80.290 168.925 80.520 175.965 ;
        RECT 80.930 168.925 81.160 175.965 ;
        RECT 81.570 168.925 81.800 175.965 ;
        RECT 82.200 175.900 82.440 175.965 ;
        RECT 82.210 168.925 82.440 175.900 ;
        RECT 75.200 168.750 75.400 168.925 ;
        RECT 76.450 168.750 76.650 168.925 ;
        RECT 77.750 168.750 77.950 168.925 ;
        RECT 79.000 168.750 79.200 168.925 ;
        RECT 80.300 168.750 80.500 168.925 ;
        RECT 81.600 168.750 81.800 168.925 ;
        RECT 72.800 167.750 81.800 168.750 ;
        RECT 85.100 167.700 87.100 176.150 ;
        RECT 75.450 167.200 75.760 167.240 ;
        RECT 76.090 167.200 76.400 167.240 ;
        RECT 76.730 167.200 77.040 167.240 ;
        RECT 77.370 167.200 77.680 167.240 ;
        RECT 78.010 167.200 78.320 167.240 ;
        RECT 78.650 167.200 78.960 167.240 ;
        RECT 79.290 167.200 79.600 167.240 ;
        RECT 79.930 167.200 80.240 167.240 ;
        RECT 80.570 167.200 80.880 167.240 ;
        RECT 81.210 167.200 81.520 167.240 ;
        RECT 81.850 167.200 82.160 167.240 ;
        RECT 82.550 167.200 82.950 167.450 ;
        RECT 75.450 167.050 82.950 167.200 ;
        RECT 85.100 167.150 87.650 167.700 ;
        RECT 75.450 167.010 82.160 167.050 ;
        RECT 75.500 167.000 82.100 167.010 ;
        RECT 60.730 165.550 72.500 165.600 ;
        RECT 58.550 165.450 72.500 165.550 ;
        RECT 58.550 165.400 61.980 165.450 ;
        RECT 52.500 159.900 52.950 160.050 ;
        RECT 31.600 158.900 32.000 159.300 ;
        RECT 30.300 131.650 30.610 131.690 ;
        RECT 23.450 131.500 30.610 131.650 ;
        RECT 23.450 131.460 24.410 131.500 ;
        RECT 24.740 131.460 25.700 131.500 ;
        RECT 26.030 131.460 26.990 131.500 ;
        RECT 30.300 131.460 30.610 131.500 ;
        RECT 23.465 131.150 26.975 131.180 ;
        RECT 29.830 131.150 31.080 131.180 ;
        RECT 31.250 131.150 31.400 137.845 ;
        RECT 32.000 133.700 32.400 133.950 ;
        RECT 34.500 133.700 34.650 159.750 ;
        RECT 52.200 159.600 52.650 159.750 ;
        RECT 51.950 159.350 52.350 159.450 ;
        RECT 35.550 159.200 52.350 159.350 ;
        RECT 35.550 158.300 35.750 159.200 ;
        RECT 51.950 159.050 52.350 159.200 ;
        RECT 52.500 158.850 52.650 159.600 ;
        RECT 47.055 158.700 49.805 158.760 ;
        RECT 52.200 158.700 52.650 158.850 ;
        RECT 45.650 158.550 51.250 158.700 ;
        RECT 35.550 157.600 35.700 158.300 ;
        RECT 35.930 158.260 39.730 158.490 ;
        RECT 39.900 158.000 40.300 158.150 ;
        RECT 39.750 157.980 40.300 158.000 ;
        RECT 35.850 157.750 40.300 157.980 ;
        RECT 35.550 156.410 35.750 157.600 ;
        RECT 35.550 156.350 35.800 156.410 ;
        RECT 35.000 142.515 35.230 155.575 ;
        RECT 35.570 150.850 35.800 156.350 ;
        RECT 35.550 150.770 35.800 150.850 ;
        RECT 39.860 151.000 40.090 156.410 ;
        RECT 40.430 151.000 40.660 155.575 ;
        RECT 39.860 150.850 40.660 151.000 ;
        RECT 39.860 150.770 40.090 150.850 ;
        RECT 35.550 147.320 35.700 150.770 ;
        RECT 35.850 149.400 39.810 149.430 ;
        RECT 35.850 149.250 39.850 149.400 ;
        RECT 35.850 149.200 40.250 149.250 ;
        RECT 39.700 148.890 40.250 149.200 ;
        RECT 35.850 148.850 40.250 148.890 ;
        RECT 35.850 148.700 39.850 148.850 ;
        RECT 35.850 148.660 39.810 148.700 ;
        RECT 35.550 147.250 35.800 147.320 ;
        RECT 35.570 141.680 35.800 147.250 ;
        RECT 39.860 141.900 40.090 147.320 ;
        RECT 40.430 142.515 40.660 150.850 ;
        RECT 45.650 148.320 45.800 158.550 ;
        RECT 47.055 158.530 49.805 158.550 ;
        RECT 46.450 158.020 50.410 158.250 ;
        RECT 46.170 155.700 46.400 157.140 ;
        RECT 46.150 155.580 46.400 155.700 ;
        RECT 46.150 153.050 46.300 155.580 ;
        RECT 46.600 154.700 46.750 158.020 ;
        RECT 50.460 155.700 50.690 157.140 ;
        RECT 50.460 155.580 50.700 155.700 ;
        RECT 46.450 154.470 50.410 154.700 ;
        RECT 46.600 154.160 46.750 154.470 ;
        RECT 46.450 153.930 50.410 154.160 ;
        RECT 46.150 152.950 46.400 153.050 ;
        RECT 46.170 151.600 46.400 152.950 ;
        RECT 46.150 151.490 46.400 151.600 ;
        RECT 46.150 148.960 46.300 151.490 ;
        RECT 46.600 150.610 46.750 153.930 ;
        RECT 50.550 153.050 50.700 155.580 ;
        RECT 50.460 151.490 50.700 153.050 ;
        RECT 46.450 150.380 50.410 150.610 ;
        RECT 46.600 150.070 46.750 150.380 ;
        RECT 46.450 149.840 50.410 150.070 ;
        RECT 46.150 148.850 46.400 148.960 ;
        RECT 40.450 141.900 40.600 142.515 ;
        RECT 39.860 141.750 40.600 141.900 ;
        RECT 39.860 141.680 40.090 141.750 ;
        RECT 39.900 140.350 40.300 140.400 ;
        RECT 39.750 140.340 40.300 140.350 ;
        RECT 35.850 140.110 40.300 140.340 ;
        RECT 39.750 140.100 40.300 140.110 ;
        RECT 39.900 140.000 40.300 140.100 ;
        RECT 35.930 139.800 39.730 139.830 ;
        RECT 40.450 139.800 40.600 141.750 ;
        RECT 45.600 139.800 45.830 148.320 ;
        RECT 46.170 147.500 46.400 148.850 ;
        RECT 46.150 147.400 46.400 147.500 ;
        RECT 46.150 144.870 46.300 147.400 ;
        RECT 46.600 146.520 46.750 149.840 ;
        RECT 50.550 148.960 50.700 151.490 ;
        RECT 50.460 147.400 50.700 148.960 ;
        RECT 51.100 148.320 51.250 158.550 ;
        RECT 46.450 146.290 50.410 146.520 ;
        RECT 46.600 145.980 46.750 146.290 ;
        RECT 46.450 145.750 50.410 145.980 ;
        RECT 46.150 144.750 46.400 144.870 ;
        RECT 46.170 143.450 46.400 144.750 ;
        RECT 46.150 143.310 46.400 143.450 ;
        RECT 46.150 140.780 46.300 143.310 ;
        RECT 46.600 142.430 46.750 145.750 ;
        RECT 50.550 144.870 50.700 147.400 ;
        RECT 50.460 143.310 50.700 144.870 ;
        RECT 46.450 142.200 50.410 142.430 ;
        RECT 46.600 141.890 46.750 142.200 ;
        RECT 46.450 141.660 50.410 141.890 ;
        RECT 46.150 140.700 46.400 140.780 ;
        RECT 35.930 139.650 45.830 139.800 ;
        RECT 35.930 139.600 39.730 139.650 ;
        RECT 35.930 138.320 39.730 138.550 ;
        RECT 39.900 138.050 40.300 138.200 ;
        RECT 39.750 138.040 40.300 138.050 ;
        RECT 35.850 137.810 40.300 138.040 ;
        RECT 39.750 137.800 40.300 137.810 ;
        RECT 32.000 133.550 34.650 133.700 ;
        RECT 13.015 131.000 16.525 131.030 ;
        RECT 19.380 131.000 20.630 131.030 ;
        RECT 20.800 131.000 31.400 131.150 ;
        RECT 31.650 133.200 34.150 133.350 ;
        RECT 12.200 130.850 20.950 131.000 ;
        RECT 23.465 130.950 26.975 131.000 ;
        RECT 29.830 130.950 31.080 131.000 ;
        RECT 12.200 127.325 12.350 130.850 ;
        RECT 13.015 130.800 16.525 130.850 ;
        RECT 19.380 130.800 20.630 130.850 ;
        RECT 17.550 130.300 17.950 130.700 ;
        RECT 13.015 128.960 16.525 129.190 ;
        RECT 13.000 128.650 13.960 128.680 ;
        RECT 14.290 128.650 15.250 128.680 ;
        RECT 15.580 128.650 16.540 128.680 ;
        RECT 17.550 128.650 17.700 130.300 ;
        RECT 19.380 128.960 20.630 129.190 ;
        RECT 23.465 129.110 26.975 129.340 ;
        RECT 29.830 129.110 31.080 129.340 ;
        RECT 31.650 129.300 31.800 133.200 ;
        RECT 32.000 132.650 32.400 132.900 ;
        RECT 32.580 132.820 33.830 133.050 ;
        RECT 34.000 132.650 34.150 133.200 ;
        RECT 32.000 132.500 32.850 132.650 ;
        RECT 33.000 132.500 34.150 132.650 ;
        RECT 32.200 129.475 32.430 132.325 ;
        RECT 32.700 131.795 32.850 132.500 ;
        RECT 33.050 132.310 33.360 132.500 ;
        RECT 32.700 131.600 33.000 131.795 ;
        RECT 32.770 130.005 33.000 131.600 ;
        RECT 33.410 130.200 33.640 131.795 ;
        RECT 33.410 130.005 33.700 130.200 ;
        RECT 33.050 129.300 33.360 129.490 ;
        RECT 31.650 129.260 33.360 129.300 ;
        RECT 33.550 129.300 33.700 130.005 ;
        RECT 33.980 129.475 34.210 132.325 ;
        RECT 35.000 130.300 35.230 137.000 ;
        RECT 35.570 130.900 35.800 136.470 ;
        RECT 35.550 130.830 35.800 130.900 ;
        RECT 39.860 131.050 40.090 136.470 ;
        RECT 40.430 131.050 40.660 137.000 ;
        RECT 39.860 130.900 40.660 131.050 ;
        RECT 39.860 130.830 40.090 130.900 ;
        RECT 35.550 129.300 35.700 130.830 ;
        RECT 40.430 130.300 40.660 130.900 ;
        RECT 39.750 129.490 40.300 129.500 ;
        RECT 31.650 129.150 33.300 129.260 ;
        RECT 33.550 129.150 35.700 129.300 ;
        RECT 35.850 129.260 40.300 129.490 ;
        RECT 39.750 129.250 40.300 129.260 ;
        RECT 23.450 128.800 24.410 128.830 ;
        RECT 24.740 128.800 25.700 128.830 ;
        RECT 26.030 128.800 26.990 128.830 ;
        RECT 30.300 128.800 30.610 128.830 ;
        RECT 19.850 128.650 20.160 128.680 ;
        RECT 21.150 128.650 30.610 128.800 ;
        RECT 13.000 128.500 21.300 128.650 ;
        RECT 23.450 128.600 24.410 128.650 ;
        RECT 24.740 128.600 25.700 128.650 ;
        RECT 26.030 128.600 26.990 128.650 ;
        RECT 13.000 128.450 13.960 128.500 ;
        RECT 14.290 128.450 15.250 128.500 ;
        RECT 15.580 128.450 16.540 128.500 ;
        RECT 17.550 128.200 17.700 128.500 ;
        RECT 19.850 128.450 20.160 128.500 ;
        RECT 17.550 127.800 17.950 128.200 ;
        RECT 21.150 127.650 21.300 128.500 ;
        RECT 27.600 127.800 28.000 128.050 ;
        RECT 14.050 127.500 19.750 127.650 ;
        RECT 12.150 119.165 12.380 127.325 ;
        RECT 14.050 126.765 14.200 127.500 ;
        RECT 16.600 126.765 16.750 127.500 ;
        RECT 12.720 119.725 12.950 126.765 ;
        RECT 14.010 119.725 14.240 126.765 ;
        RECT 15.300 119.725 15.530 126.765 ;
        RECT 16.590 119.725 16.820 126.765 ;
        RECT 12.200 119.000 12.350 119.165 ;
        RECT 12.750 119.000 12.900 119.725 ;
        RECT 15.350 119.000 15.500 119.725 ;
        RECT 17.160 119.165 17.390 127.325 ;
        RECT 17.550 126.950 17.950 127.350 ;
        RECT 12.200 118.850 15.500 119.000 ;
        RECT 12.200 117.500 12.350 118.850 ;
        RECT 13.000 118.000 13.960 118.040 ;
        RECT 14.290 118.000 15.250 118.040 ;
        RECT 15.580 118.000 16.540 118.040 ;
        RECT 17.550 118.000 17.700 126.950 ;
        RECT 19.000 119.165 19.230 127.325 ;
        RECT 19.600 126.765 19.750 127.500 ;
        RECT 20.250 127.500 21.300 127.650 ;
        RECT 20.250 126.765 20.400 127.500 ;
        RECT 19.570 119.725 19.800 126.765 ;
        RECT 20.210 119.725 20.440 126.765 ;
        RECT 20.780 119.165 21.010 127.325 ;
        RECT 20.800 118.100 20.950 119.165 ;
        RECT 19.850 118.000 20.160 118.040 ;
        RECT 12.900 117.850 20.160 118.000 ;
        RECT 13.000 117.810 13.960 117.850 ;
        RECT 14.290 117.810 15.250 117.850 ;
        RECT 15.580 117.810 16.540 117.850 ;
        RECT 19.850 117.810 20.160 117.850 ;
        RECT 20.550 117.700 20.950 118.100 ;
        RECT 13.015 117.500 16.525 117.530 ;
        RECT 19.380 117.500 20.630 117.530 ;
        RECT 20.800 117.500 20.950 117.700 ;
        RECT 12.200 117.350 20.950 117.500 ;
        RECT 12.350 117.000 12.500 117.350 ;
        RECT 13.015 117.300 16.525 117.350 ;
        RECT 19.380 117.300 20.630 117.350 ;
        RECT 21.150 117.300 21.300 127.500 ;
        RECT 24.500 127.650 28.000 127.800 ;
        RECT 22.600 119.315 22.830 127.475 ;
        RECT 24.500 126.915 24.650 127.650 ;
        RECT 27.100 126.915 27.250 127.650 ;
        RECT 23.170 119.875 23.400 126.915 ;
        RECT 24.460 119.875 24.690 126.915 ;
        RECT 25.750 119.875 25.980 126.915 ;
        RECT 27.040 119.875 27.270 126.915 ;
        RECT 22.650 119.150 22.800 119.315 ;
        RECT 23.200 119.150 23.350 119.875 ;
        RECT 25.800 119.150 25.950 119.875 ;
        RECT 27.610 119.315 27.840 127.475 ;
        RECT 22.650 119.000 25.950 119.150 ;
        RECT 22.650 117.900 22.800 119.000 ;
        RECT 23.450 118.150 24.410 118.190 ;
        RECT 24.740 118.150 25.700 118.190 ;
        RECT 26.030 118.150 26.990 118.190 ;
        RECT 28.150 118.150 28.300 128.650 ;
        RECT 30.300 128.600 30.610 128.650 ;
        RECT 29.450 127.800 29.850 128.050 ;
        RECT 31.650 127.800 31.800 129.150 ;
        RECT 39.900 129.100 40.300 129.250 ;
        RECT 32.580 128.950 33.830 128.980 ;
        RECT 35.930 128.950 39.730 128.980 ;
        RECT 40.450 128.950 40.600 130.300 ;
        RECT 45.600 128.950 45.830 139.650 ;
        RECT 46.170 139.350 46.400 140.700 ;
        RECT 46.150 139.220 46.400 139.350 ;
        RECT 46.150 136.690 46.300 139.220 ;
        RECT 46.600 138.340 46.750 141.660 ;
        RECT 50.550 140.780 50.700 143.310 ;
        RECT 50.460 139.220 50.700 140.780 ;
        RECT 46.450 138.110 50.410 138.340 ;
        RECT 46.600 137.800 46.750 138.110 ;
        RECT 46.450 137.570 50.410 137.800 ;
        RECT 46.150 136.600 46.400 136.690 ;
        RECT 46.170 135.250 46.400 136.600 ;
        RECT 46.150 135.130 46.400 135.250 ;
        RECT 46.150 132.600 46.300 135.130 ;
        RECT 46.600 134.250 46.750 137.570 ;
        RECT 50.550 136.690 50.700 139.220 ;
        RECT 50.460 135.130 50.700 136.690 ;
        RECT 46.450 134.020 50.410 134.250 ;
        RECT 46.600 133.710 46.750 134.020 ;
        RECT 46.450 133.480 50.410 133.710 ;
        RECT 46.150 132.500 46.400 132.600 ;
        RECT 46.170 131.100 46.400 132.500 ;
        RECT 32.580 128.800 45.830 128.950 ;
        RECT 32.580 128.750 33.830 128.800 ;
        RECT 35.930 128.750 39.730 128.800 ;
        RECT 29.450 127.650 30.200 127.800 ;
        RECT 29.450 119.315 29.680 127.475 ;
        RECT 30.050 126.915 30.200 127.650 ;
        RECT 30.700 127.650 31.800 127.800 ;
        RECT 30.700 126.915 30.850 127.650 ;
        RECT 30.020 119.875 30.250 126.915 ;
        RECT 30.660 119.875 30.890 126.915 ;
        RECT 31.230 119.315 31.460 127.475 ;
        RECT 31.650 121.800 31.800 127.650 ;
        RECT 35.935 127.475 39.735 127.705 ;
        RECT 45.600 127.590 45.830 128.800 ;
        RECT 46.150 131.040 46.400 131.100 ;
        RECT 46.150 128.510 46.300 131.040 ;
        RECT 46.600 130.160 46.750 133.480 ;
        RECT 50.550 132.600 50.700 135.130 ;
        RECT 50.460 131.040 50.700 132.600 ;
        RECT 46.450 129.930 50.410 130.160 ;
        RECT 46.600 129.620 46.750 129.930 ;
        RECT 46.450 129.390 50.410 129.620 ;
        RECT 46.150 128.450 46.400 128.510 ;
        RECT 39.900 127.200 40.300 127.350 ;
        RECT 39.750 127.195 40.300 127.200 ;
        RECT 35.855 127.150 40.300 127.195 ;
        RECT 35.550 127.000 40.300 127.150 ;
        RECT 32.580 121.970 33.830 122.200 ;
        RECT 31.650 121.650 32.900 121.800 ;
        RECT 33.050 121.650 33.360 121.690 ;
        RECT 32.750 121.500 33.360 121.650 ;
        RECT 30.300 118.150 30.610 118.190 ;
        RECT 23.450 118.000 30.610 118.150 ;
        RECT 23.450 117.960 24.410 118.000 ;
        RECT 24.740 117.960 25.700 118.000 ;
        RECT 26.030 117.960 26.990 118.000 ;
        RECT 30.300 117.960 30.610 118.000 ;
        RECT 22.650 117.650 23.050 117.900 ;
        RECT 23.465 117.650 26.975 117.680 ;
        RECT 29.830 117.650 31.080 117.680 ;
        RECT 31.250 117.650 31.400 119.315 ;
        RECT 32.200 118.625 32.430 121.475 ;
        RECT 32.750 120.945 32.900 121.500 ;
        RECT 33.050 121.460 33.360 121.500 ;
        RECT 32.750 120.550 33.000 120.945 ;
        RECT 32.770 119.250 33.000 120.550 ;
        RECT 32.750 119.155 33.000 119.250 ;
        RECT 33.410 119.350 33.640 120.945 ;
        RECT 33.410 119.155 33.700 119.350 ;
        RECT 32.750 118.600 32.900 119.155 ;
        RECT 33.050 118.600 33.360 118.640 ;
        RECT 32.750 118.450 33.360 118.600 ;
        RECT 33.050 118.410 33.360 118.450 ;
        RECT 33.550 118.450 33.700 119.155 ;
        RECT 33.980 118.625 34.210 121.475 ;
        RECT 35.005 119.455 35.235 126.155 ;
        RECT 35.550 125.625 35.700 127.000 ;
        RECT 35.855 126.965 40.300 127.000 ;
        RECT 39.750 126.950 40.300 126.965 ;
        RECT 35.550 125.500 35.805 125.625 ;
        RECT 35.575 120.100 35.805 125.500 ;
        RECT 35.550 119.985 35.805 120.100 ;
        RECT 39.865 120.200 40.095 125.625 ;
        RECT 40.435 120.200 40.665 126.155 ;
        RECT 39.865 120.050 40.665 120.200 ;
        RECT 39.865 119.985 40.095 120.050 ;
        RECT 35.550 118.450 35.700 119.985 ;
        RECT 40.435 119.455 40.665 120.050 ;
        RECT 35.855 118.450 39.815 118.645 ;
        RECT 33.550 118.415 39.815 118.450 ;
        RECT 33.550 118.300 36.050 118.415 ;
        RECT 32.580 118.100 33.830 118.130 ;
        RECT 35.935 118.100 39.735 118.135 ;
        RECT 40.450 118.100 40.600 119.455 ;
        RECT 45.650 118.100 45.800 127.590 ;
        RECT 46.170 127.050 46.400 128.450 ;
        RECT 46.150 126.950 46.400 127.050 ;
        RECT 46.150 124.420 46.300 126.950 ;
        RECT 46.600 126.070 46.750 129.390 ;
        RECT 50.550 128.510 50.700 131.040 ;
        RECT 50.460 128.450 50.700 128.510 ;
        RECT 51.030 135.550 51.260 148.320 ;
        RECT 52.200 135.850 52.350 158.700 ;
        RECT 52.800 145.500 52.950 159.900 ;
        RECT 58.550 149.850 58.700 165.400 ;
        RECT 60.730 165.370 61.980 165.400 ;
        RECT 64.330 165.370 65.580 165.450 ;
        RECT 67.980 165.420 69.230 165.450 ;
        RECT 68.450 165.100 68.760 165.140 ;
        RECT 61.200 165.050 61.510 165.090 ;
        RECT 64.800 165.050 65.110 165.090 ;
        RECT 60.050 164.900 65.110 165.050 ;
        RECT 60.050 162.000 60.200 164.900 ;
        RECT 61.200 164.860 61.510 164.900 ;
        RECT 64.500 163.690 64.650 164.900 ;
        RECT 64.800 164.860 65.110 164.900 ;
        RECT 68.150 164.910 68.760 165.100 ;
        RECT 68.150 164.900 68.700 164.910 ;
        RECT 68.150 163.740 68.300 164.900 ;
        RECT 68.950 163.740 69.100 165.420 ;
        RECT 60.350 163.400 60.750 163.650 ;
        RECT 60.920 163.400 61.150 163.690 ;
        RECT 60.350 163.250 61.150 163.400 ;
        RECT 60.920 163.210 61.150 163.250 ;
        RECT 61.560 163.400 61.790 163.690 ;
        RECT 61.560 163.250 62.650 163.400 ;
        RECT 61.560 163.210 61.790 163.250 ;
        RECT 61.200 162.000 61.510 162.040 ;
        RECT 60.050 161.850 61.510 162.000 ;
        RECT 61.200 161.810 61.510 161.850 ;
        RECT 62.500 159.450 62.650 163.250 ;
        RECT 64.500 163.210 64.750 163.690 ;
        RECT 65.160 163.650 65.390 163.690 ;
        RECT 68.150 163.650 68.400 163.740 ;
        RECT 65.160 163.500 68.400 163.650 ;
        RECT 65.160 163.210 65.390 163.500 ;
        RECT 68.150 163.260 68.400 163.500 ;
        RECT 68.810 163.550 69.100 163.740 ;
        RECT 70.500 164.750 72.500 165.450 ;
        RECT 73.550 165.100 73.860 165.130 ;
        RECT 74.190 165.100 74.500 165.130 ;
        RECT 74.830 165.100 75.140 165.130 ;
        RECT 75.470 165.100 75.780 165.130 ;
        RECT 76.110 165.100 76.420 165.130 ;
        RECT 76.750 165.100 77.060 165.130 ;
        RECT 77.390 165.100 77.700 165.130 ;
        RECT 78.030 165.100 78.340 165.130 ;
        RECT 78.670 165.100 78.980 165.130 ;
        RECT 79.310 165.100 79.620 165.130 ;
        RECT 79.950 165.100 80.260 165.130 ;
        RECT 80.590 165.100 80.900 165.130 ;
        RECT 81.230 165.100 81.540 165.130 ;
        RECT 81.870 165.100 82.180 165.130 ;
        RECT 82.510 165.100 82.820 165.130 ;
        RECT 83.150 165.100 83.460 165.130 ;
        RECT 83.790 165.100 84.100 165.130 ;
        RECT 73.550 164.950 84.900 165.100 ;
        RECT 73.550 164.900 73.860 164.950 ;
        RECT 74.190 164.900 74.500 164.950 ;
        RECT 74.830 164.900 75.140 164.950 ;
        RECT 75.470 164.900 75.780 164.950 ;
        RECT 76.110 164.900 76.420 164.950 ;
        RECT 76.750 164.900 77.060 164.950 ;
        RECT 77.390 164.900 77.700 164.950 ;
        RECT 78.030 164.900 78.340 164.950 ;
        RECT 78.670 164.900 78.980 164.950 ;
        RECT 79.310 164.900 79.620 164.950 ;
        RECT 79.950 164.900 80.260 164.950 ;
        RECT 80.590 164.900 80.900 164.950 ;
        RECT 81.230 164.900 81.540 164.950 ;
        RECT 81.870 164.900 82.180 164.950 ;
        RECT 82.510 164.900 82.820 164.950 ;
        RECT 83.150 164.900 83.460 164.950 ;
        RECT 83.790 164.900 84.100 164.950 ;
        RECT 70.500 163.900 83.700 164.750 ;
        RECT 84.500 164.700 84.900 164.950 ;
        RECT 68.810 163.260 69.040 163.550 ;
        RECT 64.500 162.000 64.650 163.210 ;
        RECT 68.150 162.100 68.300 163.260 ;
        RECT 68.150 162.090 68.700 162.100 ;
        RECT 64.800 162.000 65.110 162.040 ;
        RECT 64.500 161.850 65.110 162.000 ;
        RECT 68.150 161.900 68.760 162.090 ;
        RECT 68.450 161.860 68.760 161.900 ;
        RECT 64.500 160.150 64.650 161.850 ;
        RECT 64.800 161.810 65.110 161.850 ;
        RECT 64.500 159.750 64.900 160.150 ;
        RECT 62.250 159.050 62.650 159.450 ;
        RECT 62.500 158.450 62.650 159.050 ;
        RECT 70.500 159.500 72.930 163.900 ;
        RECT 73.300 163.730 73.500 163.900 ;
        RECT 74.550 163.730 74.750 163.900 ;
        RECT 75.850 163.730 76.050 163.900 ;
        RECT 77.100 163.730 77.300 163.900 ;
        RECT 78.400 163.730 78.600 163.900 ;
        RECT 79.700 163.730 79.900 163.900 ;
        RECT 80.950 163.730 81.150 163.900 ;
        RECT 82.250 163.730 82.450 163.900 ;
        RECT 83.500 163.730 83.700 163.900 ;
        RECT 73.270 163.250 73.500 163.730 ;
        RECT 73.910 163.300 74.140 163.730 ;
        RECT 73.910 163.250 74.150 163.300 ;
        RECT 74.550 163.250 74.780 163.730 ;
        RECT 75.190 163.250 75.420 163.730 ;
        RECT 75.830 163.250 76.060 163.730 ;
        RECT 76.470 163.250 76.700 163.730 ;
        RECT 77.100 163.650 77.340 163.730 ;
        RECT 77.110 163.250 77.340 163.650 ;
        RECT 77.750 163.250 77.980 163.730 ;
        RECT 78.390 163.250 78.620 163.730 ;
        RECT 79.030 163.250 79.260 163.730 ;
        RECT 79.670 163.250 79.900 163.730 ;
        RECT 80.310 163.300 80.540 163.730 ;
        RECT 80.310 163.250 80.550 163.300 ;
        RECT 80.950 163.250 81.180 163.730 ;
        RECT 81.590 163.250 81.820 163.730 ;
        RECT 82.230 163.250 82.460 163.730 ;
        RECT 82.870 163.250 83.100 163.730 ;
        RECT 83.500 163.650 83.740 163.730 ;
        RECT 83.510 163.250 83.740 163.650 ;
        RECT 84.150 163.250 84.380 163.730 ;
        RECT 73.950 163.100 74.150 163.250 ;
        RECT 75.200 163.100 75.400 163.250 ;
        RECT 76.500 163.100 76.700 163.250 ;
        RECT 77.750 163.100 77.950 163.250 ;
        RECT 79.050 163.100 79.250 163.250 ;
        RECT 80.350 163.100 80.550 163.250 ;
        RECT 81.600 163.100 81.800 163.250 ;
        RECT 82.900 163.100 83.100 163.250 ;
        RECT 84.150 163.100 84.350 163.250 ;
        RECT 85.100 163.100 87.100 167.150 ;
        RECT 113.750 167.050 114.300 167.600 ;
        RECT 115.400 167.050 115.950 167.600 ;
        RECT 73.950 163.000 87.100 163.100 ;
        RECT 73.950 162.250 149.000 163.000 ;
        RECT 73.550 162.050 73.860 162.080 ;
        RECT 74.190 162.050 74.500 162.080 ;
        RECT 74.830 162.050 75.140 162.080 ;
        RECT 75.470 162.050 75.780 162.080 ;
        RECT 76.110 162.050 76.420 162.080 ;
        RECT 76.750 162.050 77.060 162.080 ;
        RECT 77.390 162.050 77.700 162.080 ;
        RECT 78.030 162.050 78.340 162.080 ;
        RECT 78.670 162.050 78.980 162.080 ;
        RECT 79.310 162.050 79.620 162.080 ;
        RECT 79.950 162.050 80.260 162.080 ;
        RECT 80.590 162.050 80.900 162.080 ;
        RECT 81.230 162.050 81.540 162.080 ;
        RECT 81.870 162.050 82.180 162.080 ;
        RECT 82.510 162.050 82.820 162.080 ;
        RECT 83.150 162.050 83.460 162.080 ;
        RECT 83.790 162.050 84.100 162.080 ;
        RECT 73.550 161.900 84.500 162.050 ;
        RECT 73.550 161.850 84.900 161.900 ;
        RECT 73.600 161.540 84.900 161.850 ;
        RECT 73.550 161.500 84.900 161.540 ;
        RECT 73.550 161.350 84.500 161.500 ;
        RECT 73.550 161.310 73.860 161.350 ;
        RECT 74.190 161.310 74.500 161.350 ;
        RECT 74.830 161.310 75.140 161.350 ;
        RECT 75.470 161.310 75.780 161.350 ;
        RECT 76.110 161.310 76.420 161.350 ;
        RECT 76.750 161.310 77.060 161.350 ;
        RECT 77.390 161.310 77.700 161.350 ;
        RECT 78.030 161.310 78.340 161.350 ;
        RECT 78.670 161.310 78.980 161.350 ;
        RECT 79.310 161.310 79.620 161.350 ;
        RECT 79.950 161.310 80.260 161.350 ;
        RECT 80.590 161.310 80.900 161.350 ;
        RECT 81.230 161.310 81.540 161.350 ;
        RECT 81.870 161.310 82.180 161.350 ;
        RECT 82.510 161.310 82.820 161.350 ;
        RECT 83.150 161.310 83.460 161.350 ;
        RECT 83.790 161.310 84.100 161.350 ;
        RECT 85.100 161.150 149.000 162.250 ;
        RECT 73.950 161.000 149.000 161.150 ;
        RECT 73.950 160.300 87.100 161.000 ;
        RECT 73.950 160.140 74.150 160.300 ;
        RECT 75.200 160.140 75.400 160.300 ;
        RECT 76.500 160.140 76.700 160.300 ;
        RECT 77.750 160.140 77.950 160.300 ;
        RECT 79.050 160.140 79.250 160.300 ;
        RECT 80.300 160.140 80.500 160.300 ;
        RECT 81.600 160.140 81.800 160.300 ;
        RECT 82.900 160.140 83.100 160.300 ;
        RECT 84.150 160.140 84.350 160.300 ;
        RECT 73.270 159.660 73.500 160.140 ;
        RECT 73.910 160.100 74.150 160.140 ;
        RECT 73.910 159.660 74.140 160.100 ;
        RECT 74.550 159.660 74.780 160.140 ;
        RECT 75.190 159.660 75.420 160.140 ;
        RECT 75.830 159.660 76.060 160.140 ;
        RECT 76.470 159.660 76.700 160.140 ;
        RECT 77.110 159.750 77.340 160.140 ;
        RECT 77.110 159.660 77.350 159.750 ;
        RECT 77.750 159.660 77.980 160.140 ;
        RECT 78.390 159.660 78.620 160.140 ;
        RECT 79.030 159.660 79.260 160.140 ;
        RECT 79.670 159.660 79.900 160.140 ;
        RECT 80.300 160.100 80.540 160.140 ;
        RECT 80.310 159.660 80.540 160.100 ;
        RECT 80.950 159.660 81.180 160.140 ;
        RECT 81.590 159.660 81.820 160.140 ;
        RECT 82.230 159.660 82.460 160.140 ;
        RECT 82.870 159.660 83.100 160.140 ;
        RECT 83.510 159.750 83.740 160.140 ;
        RECT 83.500 159.660 83.740 159.750 ;
        RECT 84.150 159.660 84.380 160.140 ;
        RECT 73.300 159.500 73.500 159.660 ;
        RECT 74.550 159.500 74.750 159.660 ;
        RECT 75.850 159.500 76.050 159.660 ;
        RECT 77.150 159.500 77.350 159.660 ;
        RECT 78.400 159.500 78.600 159.660 ;
        RECT 79.700 159.500 79.900 159.660 ;
        RECT 80.950 159.500 81.150 159.660 ;
        RECT 82.250 159.500 82.450 159.660 ;
        RECT 83.500 159.500 83.700 159.660 ;
        RECT 70.500 158.650 83.700 159.500 ;
        RECT 73.550 158.450 73.860 158.490 ;
        RECT 74.190 158.450 74.500 158.490 ;
        RECT 74.830 158.450 75.140 158.490 ;
        RECT 75.470 158.450 75.780 158.490 ;
        RECT 76.110 158.450 76.420 158.490 ;
        RECT 76.750 158.450 77.060 158.490 ;
        RECT 77.390 158.450 77.700 158.490 ;
        RECT 78.030 158.450 78.340 158.490 ;
        RECT 78.670 158.450 78.980 158.490 ;
        RECT 79.310 158.450 79.620 158.490 ;
        RECT 79.950 158.450 80.260 158.490 ;
        RECT 80.590 158.450 80.900 158.490 ;
        RECT 81.230 158.450 81.540 158.490 ;
        RECT 81.870 158.450 82.180 158.490 ;
        RECT 82.510 158.450 82.820 158.490 ;
        RECT 83.150 158.450 83.460 158.490 ;
        RECT 83.790 158.450 84.100 158.490 ;
        RECT 84.500 158.450 84.900 158.700 ;
        RECT 62.500 158.300 84.900 158.450 ;
        RECT 73.550 158.260 84.100 158.300 ;
        RECT 73.600 158.250 84.050 158.260 ;
        RECT 75.630 149.850 77.330 149.890 ;
        RECT 79.880 149.850 81.580 149.890 ;
        RECT 58.550 149.700 81.580 149.850 ;
        RECT 73.300 149.450 73.700 149.700 ;
        RECT 75.630 149.660 77.330 149.700 ;
        RECT 77.600 149.100 77.750 149.700 ;
        RECT 77.050 149.020 77.750 149.100 ;
        RECT 75.720 147.800 75.950 149.020 ;
        RECT 74.150 147.650 75.950 147.800 ;
        RECT 74.150 147.100 74.300 147.650 ;
        RECT 75.720 147.580 75.950 147.650 ;
        RECT 77.010 148.950 77.750 149.020 ;
        RECT 79.450 149.100 79.600 149.700 ;
        RECT 79.880 149.660 81.580 149.700 ;
        RECT 79.450 149.020 80.150 149.100 ;
        RECT 79.450 148.950 80.200 149.020 ;
        RECT 77.010 147.580 77.240 148.950 ;
        RECT 79.970 147.580 80.200 148.950 ;
        RECT 81.260 147.800 81.490 149.020 ;
        RECT 82.900 147.800 83.050 158.250 ;
        RECT 81.260 147.650 83.050 147.800 ;
        RECT 81.260 147.580 81.490 147.650 ;
        RECT 76.000 147.100 76.960 147.140 ;
        RECT 80.250 147.100 81.210 147.140 ;
        RECT 74.150 146.950 81.210 147.100 ;
        RECT 52.800 145.350 74.000 145.500 ;
        RECT 73.600 145.100 74.000 145.350 ;
        RECT 52.200 135.700 59.200 135.850 ;
        RECT 51.030 135.400 58.850 135.550 ;
        RECT 50.460 127.000 50.690 128.450 ;
        RECT 51.030 127.590 51.260 135.400 ;
        RECT 54.705 134.730 57.455 134.960 ;
        RECT 54.100 134.220 58.060 134.450 ;
        RECT 53.820 131.850 54.050 133.340 ;
        RECT 53.800 131.780 54.050 131.850 ;
        RECT 53.800 129.250 53.950 131.780 ;
        RECT 54.400 130.900 54.550 134.220 ;
        RECT 58.200 133.340 58.350 135.250 ;
        RECT 58.110 133.300 58.350 133.340 ;
        RECT 58.110 131.850 58.340 133.300 ;
        RECT 58.110 131.780 58.350 131.850 ;
        RECT 54.100 130.670 58.060 130.900 ;
        RECT 54.400 130.360 54.550 130.670 ;
        RECT 54.100 130.130 58.060 130.360 ;
        RECT 53.800 127.690 54.050 129.250 ;
        RECT 50.460 126.950 50.700 127.000 ;
        RECT 50.550 126.500 50.700 126.950 ;
        RECT 53.800 126.500 53.950 127.690 ;
        RECT 54.400 126.810 54.550 130.130 ;
        RECT 58.200 129.250 58.350 131.780 ;
        RECT 58.110 129.200 58.350 129.250 ;
        RECT 58.110 127.750 58.340 129.200 ;
        RECT 58.110 127.690 58.350 127.750 ;
        RECT 54.100 126.580 58.060 126.810 ;
        RECT 50.550 126.350 53.950 126.500 ;
        RECT 46.450 125.840 50.410 126.070 ;
        RECT 46.600 125.530 46.750 125.840 ;
        RECT 46.450 125.300 50.410 125.530 ;
        RECT 46.150 124.350 46.400 124.420 ;
        RECT 46.170 122.950 46.400 124.350 ;
        RECT 46.150 122.860 46.400 122.950 ;
        RECT 46.150 120.330 46.300 122.860 ;
        RECT 46.600 121.980 46.750 125.300 ;
        RECT 50.550 124.420 50.700 126.350 ;
        RECT 53.800 125.160 53.950 126.350 ;
        RECT 54.400 126.270 54.550 126.580 ;
        RECT 54.100 126.040 58.060 126.270 ;
        RECT 50.460 124.350 50.700 124.420 ;
        RECT 50.460 122.950 50.690 124.350 ;
        RECT 50.460 122.860 50.700 122.950 ;
        RECT 46.450 121.750 50.410 121.980 ;
        RECT 46.600 121.440 46.750 121.750 ;
        RECT 46.450 121.210 50.410 121.440 ;
        RECT 46.150 120.250 46.400 120.330 ;
        RECT 46.170 118.850 46.400 120.250 ;
        RECT 32.580 117.950 45.800 118.100 ;
        RECT 32.580 117.900 33.830 117.950 ;
        RECT 35.935 117.905 39.735 117.950 ;
        RECT 22.650 117.500 31.400 117.650 ;
        RECT 45.650 117.500 45.800 117.950 ;
        RECT 46.150 118.770 46.400 118.850 ;
        RECT 23.465 117.450 26.975 117.500 ;
        RECT 29.830 117.450 31.080 117.500 ;
        RECT 46.150 117.300 46.300 118.770 ;
        RECT 46.600 117.890 46.750 121.210 ;
        RECT 50.550 120.330 50.700 122.860 ;
        RECT 50.460 120.250 50.700 120.330 ;
        RECT 50.460 118.770 50.690 120.250 ;
        RECT 46.450 117.660 50.410 117.890 ;
        RECT 21.150 117.150 46.300 117.300 ;
        RECT 12.320 116.800 38.920 117.000 ;
        RECT 12.320 113.265 12.520 116.800 ;
        RECT 12.820 114.740 13.020 116.800 ;
        RECT 13.320 115.175 13.820 115.900 ;
        RECT 13.320 115.000 13.870 115.175 ;
        RECT 13.330 114.945 13.870 115.000 ;
        RECT 12.820 114.400 13.070 114.740 ;
        RECT 12.270 113.000 12.520 113.265 ;
        RECT 12.270 108.575 12.500 113.000 ;
        RECT 12.840 106.740 13.070 114.400 ;
        RECT 14.130 107.000 14.360 114.740 ;
        RECT 14.720 113.265 14.920 116.800 ;
        RECT 18.220 116.100 18.720 116.600 ;
        RECT 15.820 115.175 16.320 115.900 ;
        RECT 15.760 115.000 16.320 115.175 ;
        RECT 18.220 115.200 18.420 116.100 ;
        RECT 18.220 115.130 18.920 115.200 ;
        RECT 18.220 115.000 19.270 115.130 ;
        RECT 15.760 114.945 16.300 115.000 ;
        RECT 18.220 114.740 18.420 115.000 ;
        RECT 18.730 114.900 19.270 115.000 ;
        RECT 14.700 108.575 14.930 113.265 ;
        RECT 15.270 107.000 15.500 114.740 ;
        RECT 14.130 106.800 15.500 107.000 ;
        RECT 14.130 106.740 14.360 106.800 ;
        RECT 15.270 106.740 15.500 106.800 ;
        RECT 16.560 107.000 16.790 114.740 ;
        RECT 18.220 114.500 18.470 114.740 ;
        RECT 17.670 113.200 17.900 113.230 ;
        RECT 17.670 113.000 17.920 113.200 ;
        RECT 17.670 108.560 17.900 113.000 ;
        RECT 18.240 107.000 18.470 114.500 ;
        RECT 16.560 106.800 18.470 107.000 ;
        RECT 16.560 106.740 16.790 106.800 ;
        RECT 18.240 106.740 18.470 106.800 ;
        RECT 19.530 107.000 19.760 114.740 ;
        RECT 20.620 113.265 20.820 116.800 ;
        RECT 21.220 114.740 21.420 116.800 ;
        RECT 21.720 115.175 22.220 115.900 ;
        RECT 21.720 115.000 22.270 115.175 ;
        RECT 21.730 114.945 22.270 115.000 ;
        RECT 21.220 114.400 21.470 114.740 ;
        RECT 20.620 113.000 20.900 113.265 ;
        RECT 20.670 108.575 20.900 113.000 ;
        RECT 19.530 106.740 19.820 107.000 ;
        RECT 21.240 106.740 21.470 114.400 ;
        RECT 22.530 107.000 22.760 114.740 ;
        RECT 23.120 113.270 23.320 116.800 ;
        RECT 26.920 116.100 27.420 116.600 ;
        RECT 24.120 115.200 24.620 115.900 ;
        RECT 24.120 115.000 26.820 115.200 ;
        RECT 27.120 115.145 27.420 116.100 ;
        RECT 27.120 115.000 27.680 115.145 ;
        RECT 24.160 114.950 24.700 115.000 ;
        RECT 26.620 114.755 26.820 115.000 ;
        RECT 27.140 114.915 27.680 115.000 ;
        RECT 23.100 108.580 23.330 113.270 ;
        RECT 23.670 107.000 23.900 114.745 ;
        RECT 22.530 106.800 23.900 107.000 ;
        RECT 22.530 106.740 22.760 106.800 ;
        RECT 23.670 106.745 23.900 106.800 ;
        RECT 24.960 107.000 25.190 114.745 ;
        RECT 26.620 114.500 26.880 114.755 ;
        RECT 26.080 108.575 26.310 113.245 ;
        RECT 26.650 107.000 26.880 114.500 ;
        RECT 24.960 106.800 26.880 107.000 ;
        RECT 24.960 106.745 25.190 106.800 ;
        RECT 26.650 106.755 26.880 106.800 ;
        RECT 27.940 107.000 28.170 114.755 ;
        RECT 29.020 113.265 29.220 116.800 ;
        RECT 29.620 114.740 29.820 116.800 ;
        RECT 30.120 115.175 30.620 115.900 ;
        RECT 30.120 115.000 30.670 115.175 ;
        RECT 30.130 114.945 30.670 115.000 ;
        RECT 29.620 114.400 29.870 114.740 ;
        RECT 29.020 113.000 29.300 113.265 ;
        RECT 29.070 108.575 29.300 113.000 ;
        RECT 27.940 106.755 28.220 107.000 ;
        RECT 19.620 106.700 19.820 106.740 ;
        RECT 19.620 106.500 20.620 106.700 ;
        RECT 19.720 106.000 20.220 106.300 ;
        RECT 20.420 106.200 20.620 106.500 ;
        RECT 20.420 106.000 22.720 106.200 ;
        RECT 12.720 105.800 20.220 106.000 ;
        RECT 12.720 104.640 12.920 105.800 ;
        RECT 13.320 105.030 13.820 105.600 ;
        RECT 13.310 104.800 13.850 105.030 ;
        RECT 15.220 104.640 15.420 105.800 ;
        RECT 15.720 105.030 16.220 105.600 ;
        RECT 15.720 104.900 16.280 105.030 ;
        RECT 15.740 104.800 16.280 104.900 ;
        RECT 17.620 104.640 17.820 105.800 ;
        RECT 18.120 105.030 18.620 105.600 ;
        RECT 18.120 104.900 18.710 105.030 ;
        RECT 18.170 104.800 18.710 104.900 ;
        RECT 20.020 104.640 20.220 105.800 ;
        RECT 22.520 105.600 22.720 106.000 ;
        RECT 24.620 106.000 25.120 106.300 ;
        RECT 28.020 106.000 28.220 106.755 ;
        RECT 29.640 106.740 29.870 114.400 ;
        RECT 30.930 107.100 31.160 114.740 ;
        RECT 31.420 113.265 31.620 116.800 ;
        RECT 32.520 115.175 33.020 115.900 ;
        RECT 32.520 115.000 33.070 115.175 ;
        RECT 32.530 114.945 33.070 115.000 ;
        RECT 31.420 113.000 31.700 113.265 ;
        RECT 31.470 108.575 31.700 113.000 ;
        RECT 32.040 107.100 32.270 114.740 ;
        RECT 30.930 106.900 32.270 107.100 ;
        RECT 30.930 106.740 31.160 106.900 ;
        RECT 32.040 106.740 32.270 106.900 ;
        RECT 33.330 107.000 33.560 114.740 ;
        RECT 33.820 113.265 34.020 116.800 ;
        RECT 34.420 114.740 34.620 116.800 ;
        RECT 34.920 115.175 35.420 115.900 ;
        RECT 34.920 115.000 35.470 115.175 ;
        RECT 34.930 114.945 35.470 115.000 ;
        RECT 34.420 114.400 34.670 114.740 ;
        RECT 33.820 113.000 34.100 113.265 ;
        RECT 33.870 108.575 34.100 113.000 ;
        RECT 33.330 106.740 33.620 107.000 ;
        RECT 34.440 106.740 34.670 114.400 ;
        RECT 35.730 107.000 35.960 114.740 ;
        RECT 36.220 113.265 36.420 116.800 ;
        RECT 38.020 116.100 38.520 116.600 ;
        RECT 37.320 115.175 37.820 115.900 ;
        RECT 37.320 115.000 37.865 115.175 ;
        RECT 37.325 114.945 37.865 115.000 ;
        RECT 38.220 114.740 38.420 116.100 ;
        RECT 36.220 113.000 36.495 113.265 ;
        RECT 36.265 108.575 36.495 113.000 ;
        RECT 36.835 107.000 37.065 114.740 ;
        RECT 35.730 106.800 37.065 107.000 ;
        RECT 35.730 106.740 35.960 106.800 ;
        RECT 36.835 106.740 37.065 106.800 ;
        RECT 38.125 114.500 38.420 114.740 ;
        RECT 38.125 106.740 38.355 114.500 ;
        RECT 38.720 110.580 38.920 116.800 ;
        RECT 39.550 116.250 39.950 116.500 ;
        RECT 46.600 116.250 46.750 117.660 ;
        RECT 47.055 117.150 49.805 117.380 ;
        RECT 39.550 116.100 50.150 116.250 ;
        RECT 39.520 115.400 40.020 115.900 ;
        RECT 39.270 112.300 39.500 112.845 ;
        RECT 39.220 111.965 39.500 112.300 ;
        RECT 39.820 112.460 40.020 115.400 ;
        RECT 44.120 113.100 44.620 113.600 ;
        RECT 44.120 112.850 44.320 113.100 ;
        RECT 42.080 112.620 46.120 112.850 ;
        RECT 39.820 112.200 40.070 112.460 ;
        RECT 48.130 112.300 48.360 112.460 ;
        RECT 39.840 112.040 40.070 112.200 ;
        RECT 48.120 112.040 48.360 112.300 ;
        RECT 39.220 111.500 39.420 111.965 ;
        RECT 48.120 111.500 48.320 112.040 ;
        RECT 39.220 111.300 49.820 111.500 ;
        RECT 45.320 110.595 49.420 110.600 ;
        RECT 38.720 110.100 39.000 110.580 ;
        RECT 41.580 110.400 49.420 110.595 ;
        RECT 41.580 110.365 45.620 110.400 ;
        RECT 39.340 110.100 39.570 110.160 ;
        RECT 38.720 109.900 39.570 110.100 ;
        RECT 47.630 110.000 47.860 110.160 ;
        RECT 38.770 109.680 39.000 109.900 ;
        RECT 39.340 109.740 39.570 109.900 ;
        RECT 47.620 109.800 49.020 110.000 ;
        RECT 47.630 109.740 47.860 109.800 ;
        RECT 48.820 108.600 49.020 109.800 ;
        RECT 48.520 108.300 49.020 108.600 ;
        RECT 47.520 108.240 49.020 108.300 ;
        RECT 39.860 108.100 49.020 108.240 ;
        RECT 39.860 108.010 47.860 108.100 ;
        RECT 39.270 107.400 39.500 107.880 ;
        RECT 48.020 107.700 48.250 107.750 ;
        RECT 49.220 107.700 49.420 110.400 ;
        RECT 48.020 107.500 49.420 107.700 ;
        RECT 39.270 107.080 39.520 107.400 ;
        RECT 48.020 107.210 48.250 107.500 ;
        RECT 48.520 107.200 49.020 107.500 ;
        RECT 33.420 106.000 33.620 106.740 ;
        RECT 39.320 106.400 39.520 107.080 ;
        RECT 39.860 106.720 47.860 106.950 ;
        RECT 39.920 106.400 40.120 106.720 ;
        RECT 49.620 106.400 49.820 111.300 ;
        RECT 39.320 106.200 49.820 106.400 ;
        RECT 24.620 105.800 32.420 106.000 ;
        RECT 33.420 105.800 48.320 106.000 ;
        RECT 20.620 105.030 21.120 105.600 ;
        RECT 22.520 105.400 23.520 105.600 ;
        RECT 20.600 104.800 21.140 105.030 ;
        RECT 22.520 104.640 22.720 105.400 ;
        RECT 23.020 105.030 23.520 105.400 ;
        RECT 23.020 104.900 23.570 105.030 ;
        RECT 23.030 104.800 23.570 104.900 ;
        RECT 24.920 104.640 25.120 105.800 ;
        RECT 25.520 105.030 26.020 105.600 ;
        RECT 25.460 104.900 26.020 105.030 ;
        RECT 25.460 104.800 26.000 104.900 ;
        RECT 27.320 104.640 27.520 105.800 ;
        RECT 27.920 105.030 28.420 105.600 ;
        RECT 27.890 104.800 28.430 105.030 ;
        RECT 29.820 104.640 30.020 105.800 ;
        RECT 30.320 105.030 30.820 105.600 ;
        RECT 30.320 104.800 30.860 105.030 ;
        RECT 32.220 104.640 32.420 105.800 ;
        RECT 32.720 105.030 33.220 105.600 ;
        RECT 32.720 104.900 33.290 105.030 ;
        RECT 32.750 104.800 33.290 104.900 ;
        RECT 38.255 104.900 44.845 104.930 ;
        RECT 48.120 104.900 48.320 105.800 ;
        RECT 38.255 104.700 48.320 104.900 ;
        RECT 12.720 104.400 13.050 104.640 ;
        RECT 12.820 96.640 13.050 104.400 ;
        RECT 14.110 96.900 14.340 104.640 ;
        RECT 15.220 104.400 15.480 104.640 ;
        RECT 14.110 96.640 14.420 96.900 ;
        RECT 15.250 96.640 15.480 104.400 ;
        RECT 16.540 96.900 16.770 104.640 ;
        RECT 17.620 104.400 17.910 104.640 ;
        RECT 16.540 96.640 16.820 96.900 ;
        RECT 17.680 96.640 17.910 104.400 ;
        RECT 18.970 96.900 19.200 104.640 ;
        RECT 20.020 104.400 20.340 104.640 ;
        RECT 18.970 96.640 19.220 96.900 ;
        RECT 20.110 96.640 20.340 104.400 ;
        RECT 21.400 96.900 21.630 104.640 ;
        RECT 22.520 104.400 22.770 104.640 ;
        RECT 21.400 96.640 21.720 96.900 ;
        RECT 22.540 96.640 22.770 104.400 ;
        RECT 23.830 96.900 24.060 104.640 ;
        RECT 24.920 104.400 25.200 104.640 ;
        RECT 23.830 96.640 24.120 96.900 ;
        RECT 24.970 96.640 25.200 104.400 ;
        RECT 26.260 96.900 26.490 104.640 ;
        RECT 27.320 104.400 27.630 104.640 ;
        RECT 26.260 96.640 26.520 96.900 ;
        RECT 27.400 96.640 27.630 104.400 ;
        RECT 28.690 96.640 28.920 104.640 ;
        RECT 29.820 104.400 30.060 104.640 ;
        RECT 29.830 96.640 30.060 104.400 ;
        RECT 31.120 96.900 31.350 104.640 ;
        RECT 32.220 104.400 32.490 104.640 ;
        RECT 31.120 96.640 31.420 96.900 ;
        RECT 32.260 96.640 32.490 104.400 ;
        RECT 33.550 96.900 33.780 104.640 ;
        RECT 48.120 104.540 48.320 104.700 ;
        RECT 34.740 103.800 34.970 104.540 ;
        RECT 48.120 104.200 48.360 104.540 ;
        RECT 34.720 103.540 34.970 103.800 ;
        RECT 48.130 103.800 48.360 104.200 ;
        RECT 48.620 103.800 49.120 104.100 ;
        RECT 48.130 103.600 49.120 103.800 ;
        RECT 48.130 103.540 48.360 103.600 ;
        RECT 34.720 102.240 34.920 103.540 ;
        RECT 37.900 102.950 45.200 103.180 ;
        RECT 36.980 102.600 41.020 102.630 ;
        RECT 44.220 102.600 44.720 102.800 ;
        RECT 36.980 102.400 44.720 102.600 ;
        RECT 44.220 102.300 44.720 102.400 ;
        RECT 44.920 102.400 45.120 102.950 ;
        RECT 49.320 102.400 49.520 106.200 ;
        RECT 34.720 101.900 34.970 102.240 ;
        RECT 34.740 101.240 34.970 101.900 ;
        RECT 43.030 101.600 43.260 102.240 ;
        RECT 44.920 102.200 49.520 102.400 ;
        RECT 43.520 101.600 44.020 101.800 ;
        RECT 43.030 101.300 44.020 101.600 ;
        RECT 43.030 101.240 43.260 101.300 ;
        RECT 44.920 101.100 45.120 102.200 ;
        RECT 43.520 100.900 45.120 101.100 ;
        RECT 41.120 100.880 43.720 100.900 ;
        RECT 36.625 100.800 43.720 100.880 ;
        RECT 34.120 100.700 43.720 100.800 ;
        RECT 34.120 100.650 41.375 100.700 ;
        RECT 34.120 100.600 36.920 100.650 ;
        RECT 34.120 98.500 34.320 100.600 ;
        RECT 36.980 100.300 41.020 100.330 ;
        RECT 44.220 100.300 44.720 100.600 ;
        RECT 36.980 100.100 44.720 100.300 ;
        RECT 34.740 99.300 34.970 99.940 ;
        RECT 34.720 98.940 34.970 99.300 ;
        RECT 43.030 99.300 43.260 99.940 ;
        RECT 43.520 99.300 44.020 99.500 ;
        RECT 43.030 99.000 44.020 99.300 ;
        RECT 43.030 98.940 43.260 99.000 ;
        RECT 34.720 98.500 34.920 98.940 ;
        RECT 36.625 98.500 41.375 98.580 ;
        RECT 34.120 98.350 41.375 98.500 ;
        RECT 34.120 98.300 36.920 98.350 ;
        RECT 33.550 96.640 33.820 96.900 ;
        RECT 12.320 96.200 12.820 96.500 ;
        RECT 13.180 96.200 13.980 96.280 ;
        RECT 12.320 96.050 13.980 96.200 ;
        RECT 12.320 96.000 13.320 96.050 ;
        RECT 14.220 95.800 14.420 96.640 ;
        RECT 14.820 96.200 15.320 96.500 ;
        RECT 15.610 96.200 16.410 96.280 ;
        RECT 14.820 96.050 16.410 96.200 ;
        RECT 14.820 96.000 15.820 96.050 ;
        RECT 16.620 95.800 16.820 96.640 ;
        RECT 17.220 96.200 17.720 96.500 ;
        RECT 18.040 96.200 18.840 96.280 ;
        RECT 17.220 96.050 18.840 96.200 ;
        RECT 17.220 96.000 18.220 96.050 ;
        RECT 19.020 95.800 19.220 96.640 ;
        RECT 19.620 96.200 20.120 96.500 ;
        RECT 20.470 96.200 21.270 96.280 ;
        RECT 19.620 96.050 21.270 96.200 ;
        RECT 19.620 96.000 20.720 96.050 ;
        RECT 21.520 95.800 21.720 96.640 ;
        RECT 22.020 96.200 22.520 96.500 ;
        RECT 22.900 96.200 23.700 96.280 ;
        RECT 23.920 96.200 24.120 96.640 ;
        RECT 22.020 96.000 24.120 96.200 ;
        RECT 24.520 96.200 25.020 96.500 ;
        RECT 25.330 96.200 26.130 96.280 ;
        RECT 24.520 96.050 26.130 96.200 ;
        RECT 24.520 96.000 25.520 96.050 ;
        RECT 26.320 95.800 26.520 96.640 ;
        RECT 26.920 96.200 27.420 96.500 ;
        RECT 27.760 96.200 28.560 96.280 ;
        RECT 26.920 96.050 28.560 96.200 ;
        RECT 26.920 96.000 27.920 96.050 ;
        RECT 28.720 95.800 28.920 96.640 ;
        RECT 29.420 96.200 29.920 96.500 ;
        RECT 30.190 96.200 30.990 96.280 ;
        RECT 29.420 96.050 30.990 96.200 ;
        RECT 29.420 96.000 30.420 96.050 ;
        RECT 31.220 95.800 31.420 96.640 ;
        RECT 31.820 96.200 32.320 96.500 ;
        RECT 32.620 96.200 33.420 96.280 ;
        RECT 31.820 96.050 33.420 96.200 ;
        RECT 31.820 96.000 32.920 96.050 ;
        RECT 33.620 95.800 33.820 96.640 ;
        RECT 34.120 96.500 34.320 98.300 ;
        RECT 36.980 98.000 41.020 98.030 ;
        RECT 44.220 98.000 44.720 98.300 ;
        RECT 36.980 97.800 44.720 98.000 ;
        RECT 34.740 97.000 34.970 97.640 ;
        RECT 34.720 96.640 34.970 97.000 ;
        RECT 43.030 96.900 43.260 97.640 ;
        RECT 43.520 96.900 44.020 97.100 ;
        RECT 43.030 96.640 44.020 96.900 ;
        RECT 34.720 96.500 34.920 96.640 ;
        RECT 34.120 96.200 34.920 96.500 ;
        RECT 43.120 96.600 44.020 96.640 ;
        RECT 36.625 96.200 41.375 96.280 ;
        RECT 34.120 96.050 41.375 96.200 ;
        RECT 34.120 96.000 36.920 96.050 ;
        RECT 43.120 95.800 43.320 96.600 ;
        RECT 14.220 95.600 43.320 95.800 ;
        RECT 44.950 95.550 45.100 100.900 ;
        RECT 44.400 95.000 45.100 95.550 ;
        RECT 44.950 85.800 45.100 95.000 ;
        RECT 50.000 90.700 50.150 116.100 ;
        RECT 53.250 103.790 53.480 124.520 ;
        RECT 53.800 123.600 54.050 125.160 ;
        RECT 53.800 121.070 53.950 123.600 ;
        RECT 54.400 122.720 54.550 126.040 ;
        RECT 58.200 125.160 58.350 127.690 ;
        RECT 58.110 125.100 58.350 125.160 ;
        RECT 58.110 123.650 58.340 125.100 ;
        RECT 58.700 124.520 58.850 135.400 ;
        RECT 59.050 132.100 59.200 135.700 ;
        RECT 73.850 135.000 74.000 145.100 ;
        RECT 74.150 143.650 74.300 146.950 ;
        RECT 76.000 146.910 76.960 146.950 ;
        RECT 80.250 146.910 81.210 146.950 ;
        RECT 75.030 144.960 77.220 145.190 ;
        RECT 79.980 144.960 82.170 145.190 ;
        RECT 75.300 144.650 75.960 144.680 ;
        RECT 76.290 144.650 76.950 144.680 ;
        RECT 80.250 144.650 80.910 144.680 ;
        RECT 81.240 144.650 81.900 144.680 ;
        RECT 75.300 144.500 78.100 144.650 ;
        RECT 75.300 144.450 75.960 144.500 ;
        RECT 76.290 144.450 76.950 144.500 ;
        RECT 74.150 143.500 77.200 143.650 ;
        RECT 74.450 135.165 74.680 143.325 ;
        RECT 75.050 142.765 75.200 143.500 ;
        RECT 77.050 142.765 77.200 143.500 ;
        RECT 75.020 135.725 75.250 142.765 ;
        RECT 76.010 135.725 76.240 142.765 ;
        RECT 77.000 135.725 77.230 142.765 ;
        RECT 76.050 135.000 76.200 135.725 ;
        RECT 77.570 135.165 77.800 143.325 ;
        RECT 73.850 134.850 76.200 135.000 ;
        RECT 75.300 134.000 75.960 134.040 ;
        RECT 76.290 134.000 76.950 134.040 ;
        RECT 77.950 134.000 78.100 144.500 ;
        RECT 79.100 144.500 81.900 144.650 ;
        RECT 78.550 134.600 78.950 134.850 ;
        RECT 79.100 134.600 79.250 144.500 ;
        RECT 80.250 144.450 80.910 144.500 ;
        RECT 81.240 144.450 81.900 144.500 ;
        RECT 82.900 143.650 83.050 147.650 ;
        RECT 80.000 143.500 83.050 143.650 ;
        RECT 83.200 145.100 83.600 145.500 ;
        RECT 79.400 135.165 79.630 143.325 ;
        RECT 80.000 142.765 80.150 143.500 ;
        RECT 82.000 142.765 82.150 143.500 ;
        RECT 79.970 135.725 80.200 142.765 ;
        RECT 80.960 135.725 81.190 142.765 ;
        RECT 81.950 135.725 82.180 142.765 ;
        RECT 81.000 134.950 81.150 135.725 ;
        RECT 82.520 135.165 82.750 143.325 ;
        RECT 83.200 134.950 83.350 145.100 ;
        RECT 81.000 134.800 83.350 134.950 ;
        RECT 78.550 134.450 79.250 134.600 ;
        RECT 78.550 134.000 78.950 134.250 ;
        RECT 75.300 133.850 78.950 134.000 ;
        RECT 79.100 134.000 79.250 134.450 ;
        RECT 80.250 134.000 80.910 134.040 ;
        RECT 81.240 134.000 81.900 134.040 ;
        RECT 79.100 133.850 81.900 134.000 ;
        RECT 75.300 133.810 75.960 133.850 ;
        RECT 76.290 133.810 76.950 133.850 ;
        RECT 80.250 133.810 80.910 133.850 ;
        RECT 81.240 133.810 81.900 133.850 ;
        RECT 75.030 133.500 77.220 133.530 ;
        RECT 79.980 133.500 82.170 133.530 ;
        RECT 75.030 133.300 82.170 133.500 ;
        RECT 59.350 132.400 59.750 132.650 ;
        RECT 60.200 132.400 60.600 132.650 ;
        RECT 59.350 132.250 60.600 132.400 ;
        RECT 76.950 132.100 77.150 133.300 ;
        RECT 78.000 132.750 78.400 133.150 ;
        RECT 78.550 132.750 78.950 133.150 ;
        RECT 59.050 131.950 77.150 132.100 ;
        RECT 59.650 131.350 60.050 131.750 ;
        RECT 62.620 131.570 75.030 131.800 ;
        RECT 59.900 128.450 60.050 131.350 ;
        RECT 60.700 131.250 68.660 131.290 ;
        RECT 68.990 131.250 76.950 131.290 ;
        RECT 77.350 131.250 77.750 131.500 ;
        RECT 60.700 131.100 78.100 131.250 ;
        RECT 60.700 131.060 68.660 131.100 ;
        RECT 68.990 131.060 76.950 131.100 ;
        RECT 77.350 128.750 77.750 129.000 ;
        RECT 60.450 128.600 77.750 128.750 ;
        RECT 58.110 123.600 58.350 123.650 ;
        RECT 54.100 122.490 58.060 122.720 ;
        RECT 54.400 122.180 54.550 122.490 ;
        RECT 54.100 121.950 58.060 122.180 ;
        RECT 53.800 119.510 54.050 121.070 ;
        RECT 53.800 116.980 53.950 119.510 ;
        RECT 54.400 118.630 54.550 121.950 ;
        RECT 58.200 121.070 58.350 123.600 ;
        RECT 58.110 121.000 58.350 121.070 ;
        RECT 58.110 119.600 58.340 121.000 ;
        RECT 58.110 119.510 58.350 119.600 ;
        RECT 54.100 118.400 58.060 118.630 ;
        RECT 54.400 118.090 54.550 118.400 ;
        RECT 54.100 117.860 58.060 118.090 ;
        RECT 53.800 115.420 54.050 116.980 ;
        RECT 53.800 112.890 53.950 115.420 ;
        RECT 54.400 114.540 54.550 117.860 ;
        RECT 58.200 116.980 58.350 119.510 ;
        RECT 58.110 116.950 58.350 116.980 ;
        RECT 58.110 115.450 58.340 116.950 ;
        RECT 58.110 115.420 58.350 115.450 ;
        RECT 54.100 114.310 58.060 114.540 ;
        RECT 54.400 114.000 54.550 114.310 ;
        RECT 54.100 113.770 58.060 114.000 ;
        RECT 53.800 111.330 54.050 112.890 ;
        RECT 53.800 108.800 53.950 111.330 ;
        RECT 54.400 110.450 54.550 113.770 ;
        RECT 58.200 112.890 58.350 115.420 ;
        RECT 58.110 112.800 58.350 112.890 ;
        RECT 58.110 111.400 58.340 112.800 ;
        RECT 58.110 111.330 58.350 111.400 ;
        RECT 54.100 110.220 58.060 110.450 ;
        RECT 54.400 109.910 54.550 110.220 ;
        RECT 54.100 109.680 58.060 109.910 ;
        RECT 53.800 107.240 54.050 108.800 ;
        RECT 53.800 104.710 53.950 107.240 ;
        RECT 54.400 106.360 54.550 109.680 ;
        RECT 58.200 108.800 58.350 111.330 ;
        RECT 58.110 108.750 58.350 108.800 ;
        RECT 58.110 107.300 58.340 108.750 ;
        RECT 58.110 107.240 58.350 107.300 ;
        RECT 54.100 106.130 58.060 106.360 ;
        RECT 54.400 105.820 54.550 106.130 ;
        RECT 54.100 105.590 58.060 105.820 ;
        RECT 53.800 103.150 54.050 104.710 ;
        RECT 53.800 100.620 53.950 103.150 ;
        RECT 54.400 102.270 54.550 105.590 ;
        RECT 58.200 104.710 58.350 107.240 ;
        RECT 58.110 104.650 58.350 104.710 ;
        RECT 58.110 103.200 58.340 104.650 ;
        RECT 58.680 103.790 58.910 124.520 ;
        RECT 59.850 113.350 60.080 128.450 ;
        RECT 60.450 127.920 60.650 128.600 ;
        RECT 77.050 127.920 77.200 128.600 ;
        RECT 60.420 113.880 60.650 127.920 ;
        RECT 68.710 113.880 68.940 127.920 ;
        RECT 77.000 113.880 77.230 127.920 ;
        RECT 59.900 112.950 60.050 113.350 ;
        RECT 68.750 112.950 68.900 113.880 ;
        RECT 77.570 113.350 77.800 128.450 ;
        RECT 77.400 112.950 77.800 113.200 ;
        RECT 59.550 112.800 77.800 112.950 ;
        RECT 59.550 108.700 59.700 112.800 ;
        RECT 60.700 110.700 68.660 110.740 ;
        RECT 68.990 110.700 76.950 110.740 ;
        RECT 60.700 110.550 77.750 110.700 ;
        RECT 60.700 110.510 68.660 110.550 ;
        RECT 68.990 110.510 76.950 110.550 ;
        RECT 77.350 110.450 77.750 110.550 ;
        RECT 77.950 110.450 78.100 131.100 ;
        RECT 77.350 110.300 78.100 110.450 ;
        RECT 62.620 110.000 75.030 110.230 ;
        RECT 59.550 108.550 77.750 108.700 ;
        RECT 58.110 103.150 58.350 103.200 ;
        RECT 54.100 102.040 58.060 102.270 ;
        RECT 54.400 101.730 54.550 102.040 ;
        RECT 54.100 101.500 58.060 101.730 ;
        RECT 53.800 99.060 54.050 100.620 ;
        RECT 53.800 96.530 53.950 99.060 ;
        RECT 54.400 98.180 54.550 101.500 ;
        RECT 58.200 100.620 58.350 103.150 ;
        RECT 58.110 100.550 58.350 100.620 ;
        RECT 58.110 99.150 58.340 100.550 ;
        RECT 58.110 99.060 58.350 99.150 ;
        RECT 54.100 97.950 58.060 98.180 ;
        RECT 54.400 97.640 54.550 97.950 ;
        RECT 54.100 97.410 58.060 97.640 ;
        RECT 53.800 96.450 54.050 96.530 ;
        RECT 53.820 94.970 54.050 96.450 ;
        RECT 54.400 94.090 54.550 97.410 ;
        RECT 58.200 96.530 58.350 99.060 ;
        RECT 58.110 96.500 58.350 96.530 ;
        RECT 58.110 95.050 58.340 96.500 ;
        RECT 58.110 94.970 58.350 95.050 ;
        RECT 54.100 93.860 58.060 94.090 ;
        RECT 47.400 90.550 50.150 90.700 ;
        RECT 47.400 89.900 47.550 90.550 ;
        RECT 48.305 90.170 51.055 90.400 ;
        RECT 47.400 89.890 47.750 89.900 ;
        RECT 53.800 89.890 54.200 89.900 ;
        RECT 54.400 89.890 54.550 93.860 ;
        RECT 54.705 93.350 57.455 93.580 ;
        RECT 58.200 93.200 58.350 94.970 ;
        RECT 58.750 93.200 58.900 103.790 ;
        RECT 58.200 93.050 58.900 93.200 ;
        RECT 54.705 90.170 57.455 90.400 ;
        RECT 47.400 89.750 51.660 89.890 ;
        RECT 46.850 86.840 47.080 89.160 ;
        RECT 47.400 88.780 47.550 89.750 ;
        RECT 47.700 89.660 51.660 89.750 ;
        RECT 53.800 89.750 58.060 89.890 ;
        RECT 53.800 89.450 53.950 89.750 ;
        RECT 54.100 89.660 58.060 89.750 ;
        RECT 51.750 89.300 53.950 89.450 ;
        RECT 51.750 88.780 51.900 89.300 ;
        RECT 47.400 88.700 47.650 88.780 ;
        RECT 47.420 87.300 47.650 88.700 ;
        RECT 47.400 87.220 47.650 87.300 ;
        RECT 51.710 87.220 51.940 88.780 ;
        RECT 47.400 86.300 47.550 87.220 ;
        RECT 52.280 86.840 52.510 89.160 ;
        RECT 53.250 86.840 53.480 89.160 ;
        RECT 53.800 88.780 53.950 89.300 ;
        RECT 53.800 88.700 54.050 88.780 ;
        RECT 53.820 87.300 54.050 88.700 ;
        RECT 53.800 87.220 54.050 87.300 ;
        RECT 47.700 86.300 51.660 86.340 ;
        RECT 47.400 86.150 51.660 86.300 ;
        RECT 47.700 86.110 51.660 86.150 ;
        RECT 48.305 85.800 51.055 85.830 ;
        RECT 52.350 85.800 52.500 86.840 ;
        RECT 53.800 86.300 53.950 87.220 ;
        RECT 54.400 86.340 54.550 89.660 ;
        RECT 58.200 88.780 58.350 93.050 ;
        RECT 58.750 89.550 58.900 93.050 ;
        RECT 59.550 89.550 59.700 108.550 ;
        RECT 62.620 108.170 75.030 108.400 ;
        RECT 77.350 108.300 77.750 108.550 ;
        RECT 60.700 107.850 68.660 107.890 ;
        RECT 68.990 107.850 76.950 107.890 ;
        RECT 77.350 107.850 77.750 108.100 ;
        RECT 77.950 107.850 78.100 110.300 ;
        RECT 60.700 107.700 78.100 107.850 ;
        RECT 60.700 107.660 68.660 107.700 ;
        RECT 68.990 107.660 76.950 107.700 ;
        RECT 77.350 105.350 77.750 105.600 ;
        RECT 60.450 105.200 77.750 105.350 ;
        RECT 59.850 89.950 60.080 105.050 ;
        RECT 60.450 104.520 60.600 105.200 ;
        RECT 77.050 104.520 77.200 105.200 ;
        RECT 60.420 90.480 60.650 104.520 ;
        RECT 68.710 90.480 68.940 104.520 ;
        RECT 77.000 90.480 77.230 104.520 ;
        RECT 59.900 89.550 60.050 89.950 ;
        RECT 68.750 89.550 68.900 90.480 ;
        RECT 77.570 89.950 77.800 105.050 ;
        RECT 77.400 89.550 77.800 89.800 ;
        RECT 58.750 89.400 77.800 89.550 ;
        RECT 58.750 89.160 58.900 89.400 ;
        RECT 58.110 88.750 58.350 88.780 ;
        RECT 58.110 87.220 58.340 88.750 ;
        RECT 58.680 86.840 58.910 89.160 ;
        RECT 60.700 87.300 68.660 87.340 ;
        RECT 68.990 87.300 76.950 87.340 ;
        RECT 77.950 87.300 78.100 107.700 ;
        RECT 60.700 87.150 78.100 87.300 ;
        RECT 78.250 129.000 78.400 132.750 ;
        RECT 78.800 129.550 78.950 132.750 ;
        RECT 80.050 132.100 80.250 133.300 ;
        RECT 80.050 131.950 97.650 132.100 ;
        RECT 82.170 131.570 94.580 131.800 ;
        RECT 79.450 131.250 79.850 131.500 ;
        RECT 80.250 131.250 88.210 131.290 ;
        RECT 88.540 131.250 96.500 131.290 ;
        RECT 79.450 131.100 96.500 131.250 ;
        RECT 80.250 131.060 88.210 131.100 ;
        RECT 88.540 131.060 96.500 131.100 ;
        RECT 97.500 130.100 97.650 131.950 ;
        RECT 98.780 130.100 100.030 130.140 ;
        RECT 102.380 130.100 103.630 130.140 ;
        RECT 105.980 130.100 107.230 130.140 ;
        RECT 97.500 129.950 107.950 130.100 ;
        RECT 98.780 129.910 100.030 129.950 ;
        RECT 102.380 129.910 103.630 129.950 ;
        RECT 105.980 129.910 107.230 129.950 ;
        RECT 99.250 129.600 99.560 129.630 ;
        RECT 102.850 129.600 103.160 129.630 ;
        RECT 106.450 129.600 106.760 129.630 ;
        RECT 78.550 129.150 78.950 129.550 ;
        RECT 78.250 128.600 78.650 129.000 ;
        RECT 78.250 105.600 78.400 128.600 ;
        RECT 78.250 105.200 78.650 105.600 ;
        RECT 78.800 105.350 78.950 129.150 ;
        RECT 98.100 129.450 99.560 129.600 ;
        RECT 79.450 128.750 79.850 129.000 ;
        RECT 98.100 128.750 98.250 129.450 ;
        RECT 99.250 129.400 99.560 129.450 ;
        RECT 101.700 129.450 103.160 129.600 ;
        RECT 79.450 128.600 98.250 128.750 ;
        RECT 100.550 128.600 100.950 128.850 ;
        RECT 79.400 113.350 79.630 128.450 ;
        RECT 80.000 127.920 80.150 128.600 ;
        RECT 96.600 127.920 96.750 128.600 ;
        RECT 79.970 113.880 80.200 127.920 ;
        RECT 88.260 113.880 88.490 127.920 ;
        RECT 96.550 113.880 96.780 127.920 ;
        RECT 79.450 113.200 79.600 113.350 ;
        RECT 79.400 112.950 79.800 113.200 ;
        RECT 88.300 112.950 88.450 113.880 ;
        RECT 97.120 113.350 97.350 128.450 ;
        RECT 98.100 119.150 98.250 128.600 ;
        RECT 99.650 128.450 100.950 128.600 ;
        RECT 98.400 120.115 98.630 128.275 ;
        RECT 99.650 127.715 99.800 128.450 ;
        RECT 98.970 120.675 99.200 127.715 ;
        RECT 99.610 120.675 99.840 127.715 ;
        RECT 99.000 119.950 99.150 120.675 ;
        RECT 100.180 120.115 100.410 128.275 ;
        RECT 97.850 118.750 98.250 119.150 ;
        RECT 98.450 119.800 99.150 119.950 ;
        RECT 98.450 117.750 98.600 119.800 ;
        RECT 98.750 118.990 99.300 119.050 ;
        RECT 98.750 118.760 99.560 118.990 ;
        RECT 98.750 118.650 99.300 118.760 ;
        RECT 98.780 118.250 100.030 118.480 ;
        RECT 101.700 118.300 101.850 129.450 ;
        RECT 102.850 129.400 103.160 129.450 ;
        RECT 105.300 129.450 106.760 129.600 ;
        RECT 104.150 128.600 104.550 128.850 ;
        RECT 103.250 128.450 104.550 128.600 ;
        RECT 102.000 120.115 102.230 128.275 ;
        RECT 103.250 127.715 103.400 128.450 ;
        RECT 102.570 120.675 102.800 127.715 ;
        RECT 103.210 120.675 103.440 127.715 ;
        RECT 102.600 119.950 102.750 120.675 ;
        RECT 103.780 120.115 104.010 128.275 ;
        RECT 101.450 117.900 101.850 118.300 ;
        RECT 102.050 119.800 102.750 119.950 ;
        RECT 102.050 117.750 102.200 119.800 ;
        RECT 102.850 118.950 103.160 118.990 ;
        RECT 105.300 118.950 105.450 129.450 ;
        RECT 106.450 129.400 106.760 129.450 ;
        RECT 105.600 120.115 105.830 128.275 ;
        RECT 106.170 120.675 106.400 127.715 ;
        RECT 106.810 120.675 107.040 127.715 ;
        RECT 106.200 119.650 106.350 120.675 ;
        RECT 105.650 119.500 106.350 119.650 ;
        RECT 106.850 119.650 107.000 120.675 ;
        RECT 107.380 120.115 107.610 128.275 ;
        RECT 107.800 122.650 107.950 129.950 ;
        RECT 107.800 122.640 109.650 122.650 ;
        RECT 107.800 122.600 110.830 122.640 ;
        RECT 107.800 122.450 116.650 122.600 ;
        RECT 109.580 122.410 110.830 122.450 ;
        RECT 108.650 122.050 109.850 122.200 ;
        RECT 110.100 122.130 111.500 122.250 ;
        RECT 108.650 121.800 109.050 122.050 ;
        RECT 109.650 121.340 109.850 122.050 ;
        RECT 110.050 122.100 111.500 122.130 ;
        RECT 110.050 121.900 110.360 122.100 ;
        RECT 109.650 121.150 110.000 121.340 ;
        RECT 107.400 119.650 107.800 119.900 ;
        RECT 106.850 119.500 107.800 119.650 ;
        RECT 109.770 119.550 110.000 121.150 ;
        RECT 110.410 121.300 110.640 121.340 ;
        RECT 110.410 120.900 111.150 121.300 ;
        RECT 110.410 119.550 110.640 120.900 ;
        RECT 105.650 119.250 106.050 119.500 ;
        RECT 106.450 118.950 106.760 118.990 ;
        RECT 110.050 118.950 110.360 118.990 ;
        RECT 111.350 118.950 111.500 122.100 ;
        RECT 111.650 120.900 112.050 121.300 ;
        RECT 102.850 118.800 104.300 118.950 ;
        RECT 102.850 118.760 103.160 118.800 ;
        RECT 102.380 118.250 103.630 118.480 ;
        RECT 104.150 118.300 104.300 118.800 ;
        RECT 105.300 118.800 111.500 118.950 ;
        RECT 104.150 117.900 104.550 118.300 ;
        RECT 105.300 117.750 105.450 118.800 ;
        RECT 106.450 118.760 106.760 118.800 ;
        RECT 110.050 118.760 110.360 118.800 ;
        RECT 105.980 118.250 107.230 118.480 ;
        RECT 98.450 117.600 105.450 117.750 ;
        RECT 105.650 117.750 106.050 118.000 ;
        RECT 105.650 117.600 115.750 117.750 ;
        RECT 98.450 114.100 98.600 117.600 ;
        RECT 101.170 117.220 113.580 117.450 ;
        RECT 115.600 116.950 115.750 117.600 ;
        RECT 115.450 116.940 115.750 116.950 ;
        RECT 99.250 116.900 107.210 116.940 ;
        RECT 107.540 116.900 115.750 116.940 ;
        RECT 99.250 116.750 115.750 116.900 ;
        RECT 99.250 116.710 107.210 116.750 ;
        RECT 107.540 116.710 115.750 116.750 ;
        RECT 115.450 116.700 115.750 116.710 ;
        RECT 79.400 112.800 88.450 112.950 ;
        RECT 80.250 110.700 88.210 110.740 ;
        RECT 88.540 110.700 96.500 110.740 ;
        RECT 79.450 110.550 96.500 110.700 ;
        RECT 79.450 110.300 79.850 110.550 ;
        RECT 80.250 110.510 88.210 110.550 ;
        RECT 88.540 110.510 96.500 110.550 ;
        RECT 82.170 110.000 94.580 110.230 ;
        RECT 98.400 108.700 98.630 114.100 ;
        RECT 115.600 113.950 115.750 116.700 ;
        RECT 99.000 113.800 115.750 113.950 ;
        RECT 99.000 113.570 99.150 113.800 ;
        RECT 115.600 113.570 115.750 113.800 ;
        RECT 79.450 108.550 98.630 108.700 ;
        RECT 79.450 108.300 79.850 108.550 ;
        RECT 82.170 108.170 94.580 108.400 ;
        RECT 79.450 107.850 79.850 108.100 ;
        RECT 80.250 107.850 88.210 107.890 ;
        RECT 88.540 107.850 96.500 107.890 ;
        RECT 79.450 107.700 96.500 107.850 ;
        RECT 80.250 107.660 88.210 107.700 ;
        RECT 88.540 107.660 96.500 107.700 ;
        RECT 97.500 105.350 97.900 105.600 ;
        RECT 78.800 105.200 97.900 105.350 ;
        RECT 60.700 87.110 68.660 87.150 ;
        RECT 68.990 87.110 76.950 87.150 ;
        RECT 77.350 86.900 77.750 87.150 ;
        RECT 54.100 86.300 58.060 86.340 ;
        RECT 53.800 86.150 58.060 86.300 ;
        RECT 54.100 86.110 58.060 86.150 ;
        RECT 54.400 86.100 54.550 86.110 ;
        RECT 54.705 85.800 57.455 85.830 ;
        RECT 58.700 85.800 58.850 86.840 ;
        RECT 62.620 86.600 75.030 86.830 ;
        RECT 44.950 85.650 58.850 85.800 ;
        RECT 48.305 85.600 51.055 85.650 ;
        RECT 54.705 85.600 57.455 85.650 ;
        RECT 44.200 85.150 44.600 85.550 ;
        RECT 44.450 66.300 44.600 85.150 ;
        RECT 49.790 84.950 72.760 84.990 ;
        RECT 77.400 84.950 77.800 85.000 ;
        RECT 49.790 84.800 77.800 84.950 ;
        RECT 49.790 84.760 72.760 84.800 ;
        RECT 77.400 84.600 77.800 84.800 ;
        RECT 45.600 84.450 46.260 84.480 ;
        RECT 46.590 84.450 47.250 84.480 ;
        RECT 47.580 84.450 48.240 84.480 ;
        RECT 48.570 84.450 49.230 84.480 ;
        RECT 49.560 84.450 50.220 84.480 ;
        RECT 50.550 84.450 51.210 84.480 ;
        RECT 51.540 84.450 52.200 84.480 ;
        RECT 52.530 84.450 53.190 84.480 ;
        RECT 53.520 84.450 54.180 84.480 ;
        RECT 54.510 84.450 55.170 84.480 ;
        RECT 55.500 84.450 56.160 84.480 ;
        RECT 56.490 84.450 57.150 84.480 ;
        RECT 57.480 84.450 58.140 84.480 ;
        RECT 58.470 84.450 59.130 84.480 ;
        RECT 59.460 84.450 60.120 84.480 ;
        RECT 60.450 84.450 61.110 84.480 ;
        RECT 61.440 84.450 62.100 84.480 ;
        RECT 62.430 84.450 63.090 84.480 ;
        RECT 63.420 84.450 64.080 84.480 ;
        RECT 64.410 84.450 65.070 84.480 ;
        RECT 65.400 84.450 66.060 84.480 ;
        RECT 66.390 84.450 67.050 84.480 ;
        RECT 67.380 84.450 68.040 84.480 ;
        RECT 68.370 84.450 69.030 84.480 ;
        RECT 69.360 84.450 70.020 84.480 ;
        RECT 70.350 84.450 71.010 84.480 ;
        RECT 71.340 84.450 72.000 84.480 ;
        RECT 72.330 84.450 72.990 84.480 ;
        RECT 73.320 84.450 73.980 84.480 ;
        RECT 74.310 84.450 74.970 84.480 ;
        RECT 75.300 84.450 75.960 84.480 ;
        RECT 76.290 84.450 76.950 84.480 ;
        RECT 45.600 84.300 78.100 84.450 ;
        RECT 45.600 84.250 46.260 84.300 ;
        RECT 46.590 84.250 47.250 84.300 ;
        RECT 47.580 84.250 48.240 84.300 ;
        RECT 48.570 84.250 49.230 84.300 ;
        RECT 49.560 84.250 50.220 84.300 ;
        RECT 50.550 84.250 51.210 84.300 ;
        RECT 51.540 84.250 52.200 84.300 ;
        RECT 52.530 84.250 53.190 84.300 ;
        RECT 53.520 84.250 54.180 84.300 ;
        RECT 54.510 84.250 55.170 84.300 ;
        RECT 55.500 84.250 56.160 84.300 ;
        RECT 56.490 84.250 57.150 84.300 ;
        RECT 57.480 84.250 58.140 84.300 ;
        RECT 58.470 84.250 59.130 84.300 ;
        RECT 59.460 84.250 60.120 84.300 ;
        RECT 60.450 84.250 61.110 84.300 ;
        RECT 61.440 84.250 62.100 84.300 ;
        RECT 62.430 84.250 63.090 84.300 ;
        RECT 63.420 84.250 64.080 84.300 ;
        RECT 64.410 84.250 65.070 84.300 ;
        RECT 65.400 84.250 66.060 84.300 ;
        RECT 66.390 84.250 67.050 84.300 ;
        RECT 67.380 84.250 68.040 84.300 ;
        RECT 68.370 84.250 69.030 84.300 ;
        RECT 69.360 84.250 70.020 84.300 ;
        RECT 70.350 84.250 71.010 84.300 ;
        RECT 71.340 84.250 72.000 84.300 ;
        RECT 72.330 84.250 72.990 84.300 ;
        RECT 73.320 84.250 73.980 84.300 ;
        RECT 74.310 84.250 74.970 84.300 ;
        RECT 75.300 84.250 75.960 84.300 ;
        RECT 76.290 84.250 76.950 84.300 ;
        RECT 77.350 81.950 77.750 82.200 ;
        RECT 45.350 81.800 77.750 81.950 ;
        RECT 44.750 66.465 44.980 81.625 ;
        RECT 45.350 81.065 45.500 81.800 ;
        RECT 47.350 81.065 47.500 81.800 ;
        RECT 49.300 81.065 49.450 81.800 ;
        RECT 51.300 81.065 51.450 81.800 ;
        RECT 53.300 81.065 53.450 81.800 ;
        RECT 55.250 81.065 55.400 81.800 ;
        RECT 57.250 81.065 57.400 81.800 ;
        RECT 59.200 81.065 59.350 81.800 ;
        RECT 61.200 81.065 61.350 81.800 ;
        RECT 63.200 81.065 63.350 81.800 ;
        RECT 65.150 81.065 65.300 81.800 ;
        RECT 67.150 81.065 67.300 81.800 ;
        RECT 69.100 81.065 69.250 81.800 ;
        RECT 71.100 81.065 71.250 81.800 ;
        RECT 73.100 81.065 73.250 81.800 ;
        RECT 75.050 81.065 75.200 81.800 ;
        RECT 77.050 81.065 77.200 81.800 ;
        RECT 45.320 67.025 45.550 81.065 ;
        RECT 46.310 67.025 46.540 81.065 ;
        RECT 47.300 67.025 47.530 81.065 ;
        RECT 48.290 67.025 48.520 81.065 ;
        RECT 49.280 67.025 49.510 81.065 ;
        RECT 50.270 67.025 50.500 81.065 ;
        RECT 51.260 67.025 51.490 81.065 ;
        RECT 52.250 67.025 52.480 81.065 ;
        RECT 53.240 67.025 53.470 81.065 ;
        RECT 54.230 67.025 54.460 81.065 ;
        RECT 55.220 67.025 55.450 81.065 ;
        RECT 56.210 67.025 56.440 81.065 ;
        RECT 57.200 67.025 57.430 81.065 ;
        RECT 58.190 67.025 58.420 81.065 ;
        RECT 59.180 67.025 59.410 81.065 ;
        RECT 60.170 67.025 60.400 81.065 ;
        RECT 61.160 67.025 61.390 81.065 ;
        RECT 62.150 67.025 62.380 81.065 ;
        RECT 63.140 67.025 63.370 81.065 ;
        RECT 64.130 67.025 64.360 81.065 ;
        RECT 65.120 67.025 65.350 81.065 ;
        RECT 66.110 67.025 66.340 81.065 ;
        RECT 67.100 67.025 67.330 81.065 ;
        RECT 68.090 67.025 68.320 81.065 ;
        RECT 69.080 67.025 69.310 81.065 ;
        RECT 70.070 67.025 70.300 81.065 ;
        RECT 71.060 67.025 71.290 81.065 ;
        RECT 72.050 67.025 72.280 81.065 ;
        RECT 73.040 67.025 73.270 81.065 ;
        RECT 74.030 67.025 74.260 81.065 ;
        RECT 75.020 67.025 75.250 81.065 ;
        RECT 76.010 67.025 76.240 81.065 ;
        RECT 77.000 67.025 77.230 81.065 ;
        RECT 46.350 66.300 46.500 67.025 ;
        RECT 48.350 66.300 48.500 67.025 ;
        RECT 50.300 66.300 50.450 67.025 ;
        RECT 52.300 66.300 52.450 67.025 ;
        RECT 54.250 66.300 54.400 67.025 ;
        RECT 56.250 66.300 56.400 67.025 ;
        RECT 58.250 66.300 58.400 67.025 ;
        RECT 60.200 66.300 60.350 67.025 ;
        RECT 62.200 66.300 62.350 67.025 ;
        RECT 64.150 66.300 64.300 67.025 ;
        RECT 66.150 66.300 66.300 67.025 ;
        RECT 68.100 66.300 68.250 67.025 ;
        RECT 70.100 66.300 70.250 67.025 ;
        RECT 72.100 66.300 72.250 67.025 ;
        RECT 74.050 66.300 74.200 67.025 ;
        RECT 76.050 66.300 76.200 67.025 ;
        RECT 77.570 66.465 77.800 81.625 ;
        RECT 44.450 66.150 77.800 66.300 ;
        RECT 44.450 42.800 44.600 66.150 ;
        RECT 77.400 65.900 77.800 66.150 ;
        RECT 45.600 63.800 46.260 63.840 ;
        RECT 46.590 63.800 47.250 63.840 ;
        RECT 47.580 63.800 48.240 63.840 ;
        RECT 48.570 63.800 49.230 63.840 ;
        RECT 49.560 63.800 50.220 63.840 ;
        RECT 50.550 63.800 51.210 63.840 ;
        RECT 51.540 63.800 52.200 63.840 ;
        RECT 52.530 63.800 53.190 63.840 ;
        RECT 53.520 63.800 54.180 63.840 ;
        RECT 54.510 63.800 55.170 63.840 ;
        RECT 55.500 63.800 56.160 63.840 ;
        RECT 56.490 63.800 57.150 63.840 ;
        RECT 57.480 63.800 58.140 63.840 ;
        RECT 58.470 63.800 59.130 63.840 ;
        RECT 59.460 63.800 60.120 63.840 ;
        RECT 60.450 63.800 61.110 63.840 ;
        RECT 61.440 63.800 62.100 63.840 ;
        RECT 62.430 63.800 63.090 63.840 ;
        RECT 63.420 63.800 64.080 63.840 ;
        RECT 64.410 63.800 65.070 63.840 ;
        RECT 65.400 63.800 66.060 63.840 ;
        RECT 66.390 63.800 67.050 63.840 ;
        RECT 67.380 63.800 68.040 63.840 ;
        RECT 68.370 63.800 69.030 63.840 ;
        RECT 69.360 63.800 70.020 63.840 ;
        RECT 70.350 63.800 71.010 63.840 ;
        RECT 71.340 63.800 72.000 63.840 ;
        RECT 72.330 63.800 72.990 63.840 ;
        RECT 73.320 63.800 73.980 63.840 ;
        RECT 74.310 63.800 74.970 63.840 ;
        RECT 75.300 63.800 75.960 63.840 ;
        RECT 76.290 63.800 76.950 63.840 ;
        RECT 77.950 63.800 78.100 84.300 ;
        RECT 45.600 63.650 78.100 63.800 ;
        RECT 45.600 63.610 46.260 63.650 ;
        RECT 46.590 63.610 47.250 63.650 ;
        RECT 47.580 63.610 48.240 63.650 ;
        RECT 48.570 63.610 49.230 63.650 ;
        RECT 49.560 63.610 50.220 63.650 ;
        RECT 50.550 63.610 51.210 63.650 ;
        RECT 51.540 63.610 52.200 63.650 ;
        RECT 52.530 63.610 53.190 63.650 ;
        RECT 53.520 63.610 54.180 63.650 ;
        RECT 54.510 63.610 55.170 63.650 ;
        RECT 55.500 63.610 56.160 63.650 ;
        RECT 56.490 63.610 57.150 63.650 ;
        RECT 57.480 63.610 58.140 63.650 ;
        RECT 58.470 63.610 59.130 63.650 ;
        RECT 59.460 63.610 60.120 63.650 ;
        RECT 60.450 63.610 61.110 63.650 ;
        RECT 61.440 63.610 62.100 63.650 ;
        RECT 62.430 63.610 63.090 63.650 ;
        RECT 63.420 63.610 64.080 63.650 ;
        RECT 64.410 63.610 65.070 63.650 ;
        RECT 65.400 63.610 66.060 63.650 ;
        RECT 66.390 63.610 67.050 63.650 ;
        RECT 67.380 63.610 68.040 63.650 ;
        RECT 68.370 63.610 69.030 63.650 ;
        RECT 69.360 63.610 70.020 63.650 ;
        RECT 70.350 63.610 71.010 63.650 ;
        RECT 71.340 63.610 72.000 63.650 ;
        RECT 72.330 63.610 72.990 63.650 ;
        RECT 73.320 63.610 73.980 63.650 ;
        RECT 74.310 63.610 74.970 63.650 ;
        RECT 75.300 63.610 75.960 63.650 ;
        RECT 76.290 63.610 76.950 63.650 ;
        RECT 77.700 63.400 78.100 63.650 ;
        RECT 49.790 63.100 72.760 63.330 ;
        RECT 77.950 62.500 78.100 63.400 ;
        RECT 44.750 61.650 45.300 62.200 ;
        RECT 77.700 62.100 78.100 62.500 ;
        RECT 78.250 82.200 78.400 105.200 ;
        RECT 78.800 82.750 78.950 105.200 ;
        RECT 79.400 89.950 79.630 105.050 ;
        RECT 80.000 104.520 80.150 105.200 ;
        RECT 96.600 104.520 96.750 105.200 ;
        RECT 79.970 90.480 80.200 104.520 ;
        RECT 88.260 90.480 88.490 104.520 ;
        RECT 96.550 90.480 96.780 104.520 ;
        RECT 79.450 89.800 79.600 89.950 ;
        RECT 79.400 89.550 79.800 89.800 ;
        RECT 88.300 89.550 88.450 90.480 ;
        RECT 97.120 89.950 97.350 105.050 ;
        RECT 98.400 99.200 98.630 108.550 ;
        RECT 98.970 99.530 99.200 113.570 ;
        RECT 107.260 99.530 107.490 113.570 ;
        RECT 115.550 99.530 115.780 113.570 ;
        RECT 107.300 99.200 107.450 99.530 ;
        RECT 98.400 99.050 107.450 99.200 ;
        RECT 98.400 99.000 98.630 99.050 ;
        RECT 115.600 96.400 115.750 99.530 ;
        RECT 116.120 99.000 116.350 114.100 ;
        RECT 115.450 96.390 115.750 96.400 ;
        RECT 99.250 96.350 107.210 96.390 ;
        RECT 107.540 96.350 115.750 96.390 ;
        RECT 97.500 96.200 115.750 96.350 ;
        RECT 79.400 89.400 88.450 89.550 ;
        RECT 80.250 87.300 88.210 87.340 ;
        RECT 88.540 87.300 96.500 87.340 ;
        RECT 97.500 87.300 97.650 96.200 ;
        RECT 99.250 96.160 107.210 96.200 ;
        RECT 107.540 96.160 115.500 96.200 ;
        RECT 101.170 95.650 113.580 95.880 ;
        RECT 116.500 94.850 116.650 122.450 ;
        RECT 79.450 87.150 97.650 87.300 ;
        RECT 112.250 94.700 116.650 94.850 ;
        RECT 79.450 86.900 79.850 87.150 ;
        RECT 80.250 87.110 88.210 87.150 ;
        RECT 88.540 87.110 96.500 87.150 ;
        RECT 82.170 86.600 94.580 86.830 ;
        RECT 79.400 84.990 84.500 85.000 ;
        RECT 79.400 84.950 107.410 84.990 ;
        RECT 112.250 84.950 112.400 94.700 ;
        RECT 79.400 84.850 112.400 84.950 ;
        RECT 79.400 84.600 79.800 84.850 ;
        RECT 84.440 84.800 112.400 84.850 ;
        RECT 84.440 84.760 107.410 84.800 ;
        RECT 80.250 84.450 80.910 84.480 ;
        RECT 81.240 84.450 81.900 84.480 ;
        RECT 82.230 84.450 82.890 84.480 ;
        RECT 83.220 84.450 83.880 84.480 ;
        RECT 84.210 84.450 84.870 84.480 ;
        RECT 85.200 84.450 85.860 84.480 ;
        RECT 86.190 84.450 86.850 84.480 ;
        RECT 87.180 84.450 87.840 84.480 ;
        RECT 88.170 84.450 88.830 84.480 ;
        RECT 89.160 84.450 89.820 84.480 ;
        RECT 90.150 84.450 90.810 84.480 ;
        RECT 91.140 84.450 91.800 84.480 ;
        RECT 92.130 84.450 92.790 84.480 ;
        RECT 93.120 84.450 93.780 84.480 ;
        RECT 94.110 84.450 94.770 84.480 ;
        RECT 95.100 84.450 95.760 84.480 ;
        RECT 96.090 84.450 96.750 84.480 ;
        RECT 97.080 84.450 97.740 84.480 ;
        RECT 98.070 84.450 98.730 84.480 ;
        RECT 99.060 84.450 99.720 84.480 ;
        RECT 100.050 84.450 100.710 84.480 ;
        RECT 101.040 84.450 101.700 84.480 ;
        RECT 102.030 84.450 102.690 84.480 ;
        RECT 103.020 84.450 103.680 84.480 ;
        RECT 104.010 84.450 104.670 84.480 ;
        RECT 105.000 84.450 105.660 84.480 ;
        RECT 105.990 84.450 106.650 84.480 ;
        RECT 106.980 84.450 107.640 84.480 ;
        RECT 107.970 84.450 108.630 84.480 ;
        RECT 108.960 84.450 109.620 84.480 ;
        RECT 109.950 84.450 110.610 84.480 ;
        RECT 110.940 84.450 111.600 84.480 ;
        RECT 78.550 82.350 78.950 82.750 ;
        RECT 78.250 81.800 78.650 82.200 ;
        RECT 44.750 58.450 44.900 61.650 ;
        RECT 49.790 61.260 72.760 61.490 ;
        RECT 45.600 60.950 46.260 60.980 ;
        RECT 46.590 60.950 47.250 60.980 ;
        RECT 47.580 60.950 48.240 60.980 ;
        RECT 48.570 60.950 49.230 60.980 ;
        RECT 49.560 60.950 50.220 60.980 ;
        RECT 50.550 60.950 51.210 60.980 ;
        RECT 51.540 60.950 52.200 60.980 ;
        RECT 52.530 60.950 53.190 60.980 ;
        RECT 53.520 60.950 54.180 60.980 ;
        RECT 54.510 60.950 55.170 60.980 ;
        RECT 55.500 60.950 56.160 60.980 ;
        RECT 56.490 60.950 57.150 60.980 ;
        RECT 57.480 60.950 58.140 60.980 ;
        RECT 58.470 60.950 59.130 60.980 ;
        RECT 59.460 60.950 60.120 60.980 ;
        RECT 60.450 60.950 61.110 60.980 ;
        RECT 61.440 60.950 62.100 60.980 ;
        RECT 62.430 60.950 63.090 60.980 ;
        RECT 63.420 60.950 64.080 60.980 ;
        RECT 64.410 60.950 65.070 60.980 ;
        RECT 65.400 60.950 66.060 60.980 ;
        RECT 66.390 60.950 67.050 60.980 ;
        RECT 67.380 60.950 68.040 60.980 ;
        RECT 68.370 60.950 69.030 60.980 ;
        RECT 69.360 60.950 70.020 60.980 ;
        RECT 70.350 60.950 71.010 60.980 ;
        RECT 71.340 60.950 72.000 60.980 ;
        RECT 72.330 60.950 72.990 60.980 ;
        RECT 73.320 60.950 73.980 60.980 ;
        RECT 74.310 60.950 74.970 60.980 ;
        RECT 75.300 60.950 75.960 60.980 ;
        RECT 76.290 60.950 76.950 60.980 ;
        RECT 77.700 60.950 78.100 61.200 ;
        RECT 45.600 60.800 78.100 60.950 ;
        RECT 45.600 60.750 46.260 60.800 ;
        RECT 46.590 60.750 47.250 60.800 ;
        RECT 47.580 60.750 48.240 60.800 ;
        RECT 48.570 60.750 49.230 60.800 ;
        RECT 49.560 60.750 50.220 60.800 ;
        RECT 50.550 60.750 51.210 60.800 ;
        RECT 51.540 60.750 52.200 60.800 ;
        RECT 52.530 60.750 53.190 60.800 ;
        RECT 53.520 60.750 54.180 60.800 ;
        RECT 54.510 60.750 55.170 60.800 ;
        RECT 55.500 60.750 56.160 60.800 ;
        RECT 56.490 60.750 57.150 60.800 ;
        RECT 57.480 60.750 58.140 60.800 ;
        RECT 58.470 60.750 59.130 60.800 ;
        RECT 59.460 60.750 60.120 60.800 ;
        RECT 60.450 60.750 61.110 60.800 ;
        RECT 61.440 60.750 62.100 60.800 ;
        RECT 62.430 60.750 63.090 60.800 ;
        RECT 63.420 60.750 64.080 60.800 ;
        RECT 64.410 60.750 65.070 60.800 ;
        RECT 65.400 60.750 66.060 60.800 ;
        RECT 66.390 60.750 67.050 60.800 ;
        RECT 67.380 60.750 68.040 60.800 ;
        RECT 68.370 60.750 69.030 60.800 ;
        RECT 69.360 60.750 70.020 60.800 ;
        RECT 70.350 60.750 71.010 60.800 ;
        RECT 71.340 60.750 72.000 60.800 ;
        RECT 72.330 60.750 72.990 60.800 ;
        RECT 73.320 60.750 73.980 60.800 ;
        RECT 74.310 60.750 74.970 60.800 ;
        RECT 75.300 60.750 75.960 60.800 ;
        RECT 76.290 60.750 76.950 60.800 ;
        RECT 77.350 58.450 77.750 58.700 ;
        RECT 44.750 58.300 77.750 58.450 ;
        RECT 44.750 42.965 44.980 58.125 ;
        RECT 45.350 57.565 45.500 58.300 ;
        RECT 47.350 57.565 47.500 58.300 ;
        RECT 49.300 57.565 49.450 58.300 ;
        RECT 51.300 57.565 51.450 58.300 ;
        RECT 53.300 57.565 53.450 58.300 ;
        RECT 55.250 57.565 55.400 58.300 ;
        RECT 57.250 57.565 57.400 58.300 ;
        RECT 59.200 57.565 59.350 58.300 ;
        RECT 61.200 57.565 61.350 58.300 ;
        RECT 63.200 57.565 63.350 58.300 ;
        RECT 65.150 57.565 65.300 58.300 ;
        RECT 67.150 57.565 67.300 58.300 ;
        RECT 69.100 57.565 69.250 58.300 ;
        RECT 71.100 57.565 71.250 58.300 ;
        RECT 73.100 57.565 73.250 58.300 ;
        RECT 75.050 57.565 75.200 58.300 ;
        RECT 77.050 57.565 77.200 58.300 ;
        RECT 45.320 43.525 45.550 57.565 ;
        RECT 46.310 43.525 46.540 57.565 ;
        RECT 47.300 43.525 47.530 57.565 ;
        RECT 48.290 43.525 48.520 57.565 ;
        RECT 49.280 43.525 49.510 57.565 ;
        RECT 50.270 43.525 50.500 57.565 ;
        RECT 51.260 43.525 51.490 57.565 ;
        RECT 52.250 43.525 52.480 57.565 ;
        RECT 53.240 43.525 53.470 57.565 ;
        RECT 54.230 43.525 54.460 57.565 ;
        RECT 55.220 43.525 55.450 57.565 ;
        RECT 56.210 43.525 56.440 57.565 ;
        RECT 57.200 43.525 57.430 57.565 ;
        RECT 58.190 43.525 58.420 57.565 ;
        RECT 59.180 43.525 59.410 57.565 ;
        RECT 60.170 43.525 60.400 57.565 ;
        RECT 61.160 43.525 61.390 57.565 ;
        RECT 62.150 43.525 62.380 57.565 ;
        RECT 63.140 43.525 63.370 57.565 ;
        RECT 64.130 43.525 64.360 57.565 ;
        RECT 65.120 43.525 65.350 57.565 ;
        RECT 66.110 43.525 66.340 57.565 ;
        RECT 67.100 43.525 67.330 57.565 ;
        RECT 68.090 43.525 68.320 57.565 ;
        RECT 69.080 43.525 69.310 57.565 ;
        RECT 70.070 43.525 70.300 57.565 ;
        RECT 71.060 43.525 71.290 57.565 ;
        RECT 72.050 43.525 72.280 57.565 ;
        RECT 73.040 43.525 73.270 57.565 ;
        RECT 74.030 43.525 74.260 57.565 ;
        RECT 75.020 43.525 75.250 57.565 ;
        RECT 76.010 43.525 76.240 57.565 ;
        RECT 77.000 43.525 77.230 57.565 ;
        RECT 46.350 42.800 46.500 43.525 ;
        RECT 48.350 42.800 48.500 43.525 ;
        RECT 50.300 42.800 50.450 43.525 ;
        RECT 52.300 42.800 52.450 43.525 ;
        RECT 54.250 42.800 54.400 43.525 ;
        RECT 56.250 42.800 56.400 43.525 ;
        RECT 58.250 42.800 58.400 43.525 ;
        RECT 60.200 42.800 60.350 43.525 ;
        RECT 62.200 42.800 62.350 43.525 ;
        RECT 64.150 42.800 64.300 43.525 ;
        RECT 66.150 42.800 66.300 43.525 ;
        RECT 68.100 42.800 68.250 43.525 ;
        RECT 70.100 42.800 70.250 43.525 ;
        RECT 72.100 42.800 72.250 43.525 ;
        RECT 74.050 42.800 74.200 43.525 ;
        RECT 76.050 42.800 76.200 43.525 ;
        RECT 77.570 42.965 77.800 58.125 ;
        RECT 44.450 42.650 77.800 42.800 ;
        RECT 77.400 42.400 77.800 42.650 ;
        RECT 45.600 40.300 46.260 40.340 ;
        RECT 46.590 40.300 47.250 40.340 ;
        RECT 47.580 40.300 48.240 40.340 ;
        RECT 48.570 40.300 49.230 40.340 ;
        RECT 49.560 40.300 50.220 40.340 ;
        RECT 50.550 40.300 51.210 40.340 ;
        RECT 51.540 40.300 52.200 40.340 ;
        RECT 52.530 40.300 53.190 40.340 ;
        RECT 53.520 40.300 54.180 40.340 ;
        RECT 54.510 40.300 55.170 40.340 ;
        RECT 55.500 40.300 56.160 40.340 ;
        RECT 56.490 40.300 57.150 40.340 ;
        RECT 57.480 40.300 58.140 40.340 ;
        RECT 58.470 40.300 59.130 40.340 ;
        RECT 59.460 40.300 60.120 40.340 ;
        RECT 60.450 40.300 61.110 40.340 ;
        RECT 61.440 40.300 62.100 40.340 ;
        RECT 62.430 40.300 63.090 40.340 ;
        RECT 63.420 40.300 64.080 40.340 ;
        RECT 64.410 40.300 65.070 40.340 ;
        RECT 65.400 40.300 66.060 40.340 ;
        RECT 66.390 40.300 67.050 40.340 ;
        RECT 67.380 40.300 68.040 40.340 ;
        RECT 68.370 40.300 69.030 40.340 ;
        RECT 69.360 40.300 70.020 40.340 ;
        RECT 70.350 40.300 71.010 40.340 ;
        RECT 71.340 40.300 72.000 40.340 ;
        RECT 72.330 40.300 72.990 40.340 ;
        RECT 73.320 40.300 73.980 40.340 ;
        RECT 74.310 40.300 74.970 40.340 ;
        RECT 75.300 40.300 75.960 40.340 ;
        RECT 76.290 40.300 76.950 40.340 ;
        RECT 77.950 40.300 78.100 60.800 ;
        RECT 78.250 58.700 78.400 81.800 ;
        RECT 78.800 59.250 78.950 82.350 ;
        RECT 79.100 84.300 111.600 84.450 ;
        RECT 79.100 63.800 79.250 84.300 ;
        RECT 80.250 84.250 80.910 84.300 ;
        RECT 81.240 84.250 81.900 84.300 ;
        RECT 82.230 84.250 82.890 84.300 ;
        RECT 83.220 84.250 83.880 84.300 ;
        RECT 84.210 84.250 84.870 84.300 ;
        RECT 85.200 84.250 85.860 84.300 ;
        RECT 86.190 84.250 86.850 84.300 ;
        RECT 87.180 84.250 87.840 84.300 ;
        RECT 88.170 84.250 88.830 84.300 ;
        RECT 89.160 84.250 89.820 84.300 ;
        RECT 90.150 84.250 90.810 84.300 ;
        RECT 91.140 84.250 91.800 84.300 ;
        RECT 92.130 84.250 92.790 84.300 ;
        RECT 93.120 84.250 93.780 84.300 ;
        RECT 94.110 84.250 94.770 84.300 ;
        RECT 95.100 84.250 95.760 84.300 ;
        RECT 96.090 84.250 96.750 84.300 ;
        RECT 97.080 84.250 97.740 84.300 ;
        RECT 98.070 84.250 98.730 84.300 ;
        RECT 99.060 84.250 99.720 84.300 ;
        RECT 100.050 84.250 100.710 84.300 ;
        RECT 101.040 84.250 101.700 84.300 ;
        RECT 102.030 84.250 102.690 84.300 ;
        RECT 103.020 84.250 103.680 84.300 ;
        RECT 104.010 84.250 104.670 84.300 ;
        RECT 105.000 84.250 105.660 84.300 ;
        RECT 105.990 84.250 106.650 84.300 ;
        RECT 106.980 84.250 107.640 84.300 ;
        RECT 107.970 84.250 108.630 84.300 ;
        RECT 108.960 84.250 109.620 84.300 ;
        RECT 109.950 84.250 110.610 84.300 ;
        RECT 110.940 84.250 111.600 84.300 ;
        RECT 79.450 81.950 79.850 82.200 ;
        RECT 79.450 81.800 111.850 81.950 ;
        RECT 79.400 66.465 79.630 81.625 ;
        RECT 80.000 81.065 80.150 81.800 ;
        RECT 82.000 81.065 82.150 81.800 ;
        RECT 83.950 81.065 84.100 81.800 ;
        RECT 85.950 81.065 86.100 81.800 ;
        RECT 87.950 81.065 88.100 81.800 ;
        RECT 89.900 81.065 90.050 81.800 ;
        RECT 91.900 81.065 92.050 81.800 ;
        RECT 93.850 81.065 94.000 81.800 ;
        RECT 95.850 81.065 96.000 81.800 ;
        RECT 97.850 81.065 98.000 81.800 ;
        RECT 99.800 81.065 99.950 81.800 ;
        RECT 101.800 81.065 101.950 81.800 ;
        RECT 103.750 81.065 103.900 81.800 ;
        RECT 105.750 81.065 105.900 81.800 ;
        RECT 107.750 81.065 107.900 81.800 ;
        RECT 109.700 81.065 109.850 81.800 ;
        RECT 111.700 81.065 111.850 81.800 ;
        RECT 112.250 81.625 112.400 84.800 ;
        RECT 79.970 67.025 80.200 81.065 ;
        RECT 80.960 67.025 81.190 81.065 ;
        RECT 81.950 67.025 82.180 81.065 ;
        RECT 82.940 67.025 83.170 81.065 ;
        RECT 83.930 67.025 84.160 81.065 ;
        RECT 84.920 67.025 85.150 81.065 ;
        RECT 85.910 67.025 86.140 81.065 ;
        RECT 86.900 67.025 87.130 81.065 ;
        RECT 87.890 67.025 88.120 81.065 ;
        RECT 88.880 67.025 89.110 81.065 ;
        RECT 89.870 67.025 90.100 81.065 ;
        RECT 90.860 67.025 91.090 81.065 ;
        RECT 91.850 67.025 92.080 81.065 ;
        RECT 92.840 67.025 93.070 81.065 ;
        RECT 93.830 67.025 94.060 81.065 ;
        RECT 94.820 67.025 95.050 81.065 ;
        RECT 95.810 67.025 96.040 81.065 ;
        RECT 96.800 67.025 97.030 81.065 ;
        RECT 97.790 67.025 98.020 81.065 ;
        RECT 98.780 67.025 99.010 81.065 ;
        RECT 99.770 67.025 100.000 81.065 ;
        RECT 100.760 67.025 100.990 81.065 ;
        RECT 101.750 67.025 101.980 81.065 ;
        RECT 102.740 67.025 102.970 81.065 ;
        RECT 103.730 67.025 103.960 81.065 ;
        RECT 104.720 67.025 104.950 81.065 ;
        RECT 105.710 67.025 105.940 81.065 ;
        RECT 106.700 67.025 106.930 81.065 ;
        RECT 107.690 67.025 107.920 81.065 ;
        RECT 108.680 67.025 108.910 81.065 ;
        RECT 109.670 67.025 109.900 81.065 ;
        RECT 110.660 67.025 110.890 81.065 ;
        RECT 111.650 67.025 111.880 81.065 ;
        RECT 81.000 66.300 81.150 67.025 ;
        RECT 83.000 66.300 83.150 67.025 ;
        RECT 84.950 66.300 85.100 67.025 ;
        RECT 86.950 66.300 87.100 67.025 ;
        RECT 88.900 66.300 89.050 67.025 ;
        RECT 90.900 66.300 91.050 67.025 ;
        RECT 92.900 66.300 93.050 67.025 ;
        RECT 94.850 66.300 95.000 67.025 ;
        RECT 96.850 66.300 97.000 67.025 ;
        RECT 98.800 66.300 98.950 67.025 ;
        RECT 100.800 66.300 100.950 67.025 ;
        RECT 102.750 66.300 102.900 67.025 ;
        RECT 104.750 66.300 104.900 67.025 ;
        RECT 106.750 66.300 106.900 67.025 ;
        RECT 108.700 66.300 108.850 67.025 ;
        RECT 110.700 66.300 110.850 67.025 ;
        RECT 112.220 66.465 112.450 81.625 ;
        RECT 79.400 66.150 110.850 66.300 ;
        RECT 79.400 65.900 79.800 66.150 ;
        RECT 80.250 63.800 80.910 63.840 ;
        RECT 81.240 63.800 81.900 63.840 ;
        RECT 82.230 63.800 82.890 63.840 ;
        RECT 83.220 63.800 83.880 63.840 ;
        RECT 84.210 63.800 84.870 63.840 ;
        RECT 85.200 63.800 85.860 63.840 ;
        RECT 86.190 63.800 86.850 63.840 ;
        RECT 87.180 63.800 87.840 63.840 ;
        RECT 88.170 63.800 88.830 63.840 ;
        RECT 89.160 63.800 89.820 63.840 ;
        RECT 90.150 63.800 90.810 63.840 ;
        RECT 91.140 63.800 91.800 63.840 ;
        RECT 92.130 63.800 92.790 63.840 ;
        RECT 93.120 63.800 93.780 63.840 ;
        RECT 94.110 63.800 94.770 63.840 ;
        RECT 95.100 63.800 95.760 63.840 ;
        RECT 96.090 63.800 96.750 63.840 ;
        RECT 97.080 63.800 97.740 63.840 ;
        RECT 98.070 63.800 98.730 63.840 ;
        RECT 99.060 63.800 99.720 63.840 ;
        RECT 100.050 63.800 100.710 63.840 ;
        RECT 101.040 63.800 101.700 63.840 ;
        RECT 102.030 63.800 102.690 63.840 ;
        RECT 103.020 63.800 103.680 63.840 ;
        RECT 104.010 63.800 104.670 63.840 ;
        RECT 105.000 63.800 105.660 63.840 ;
        RECT 105.990 63.800 106.650 63.840 ;
        RECT 106.980 63.800 107.640 63.840 ;
        RECT 107.970 63.800 108.630 63.840 ;
        RECT 108.960 63.800 109.620 63.840 ;
        RECT 109.950 63.800 110.610 63.840 ;
        RECT 110.940 63.800 111.600 63.840 ;
        RECT 79.100 63.650 111.600 63.800 ;
        RECT 79.100 63.400 79.500 63.650 ;
        RECT 80.250 63.610 80.910 63.650 ;
        RECT 81.240 63.610 81.900 63.650 ;
        RECT 82.230 63.610 82.890 63.650 ;
        RECT 83.220 63.610 83.880 63.650 ;
        RECT 84.210 63.610 84.870 63.650 ;
        RECT 85.200 63.610 85.860 63.650 ;
        RECT 86.190 63.610 86.850 63.650 ;
        RECT 87.180 63.610 87.840 63.650 ;
        RECT 88.170 63.610 88.830 63.650 ;
        RECT 89.160 63.610 89.820 63.650 ;
        RECT 90.150 63.610 90.810 63.650 ;
        RECT 91.140 63.610 91.800 63.650 ;
        RECT 92.130 63.610 92.790 63.650 ;
        RECT 93.120 63.610 93.780 63.650 ;
        RECT 94.110 63.610 94.770 63.650 ;
        RECT 95.100 63.610 95.760 63.650 ;
        RECT 96.090 63.610 96.750 63.650 ;
        RECT 97.080 63.610 97.740 63.650 ;
        RECT 98.070 63.610 98.730 63.650 ;
        RECT 99.060 63.610 99.720 63.650 ;
        RECT 100.050 63.610 100.710 63.650 ;
        RECT 101.040 63.610 101.700 63.650 ;
        RECT 102.030 63.610 102.690 63.650 ;
        RECT 103.020 63.610 103.680 63.650 ;
        RECT 104.010 63.610 104.670 63.650 ;
        RECT 105.000 63.610 105.660 63.650 ;
        RECT 105.990 63.610 106.650 63.650 ;
        RECT 106.980 63.610 107.640 63.650 ;
        RECT 107.970 63.610 108.630 63.650 ;
        RECT 108.960 63.610 109.620 63.650 ;
        RECT 109.950 63.610 110.610 63.650 ;
        RECT 110.940 63.610 111.600 63.650 ;
        RECT 84.440 63.300 107.410 63.330 ;
        RECT 112.250 63.300 112.400 66.465 ;
        RECT 84.440 63.150 112.400 63.300 ;
        RECT 84.440 63.100 107.410 63.150 ;
        RECT 84.440 61.450 107.410 61.490 ;
        RECT 112.250 61.450 112.400 63.150 ;
        RECT 84.440 61.300 112.400 61.450 ;
        RECT 84.440 61.260 107.410 61.300 ;
        RECT 78.550 58.850 78.950 59.250 ;
        RECT 79.100 60.950 79.500 61.200 ;
        RECT 80.250 60.950 80.910 60.980 ;
        RECT 81.240 60.950 81.900 60.980 ;
        RECT 82.230 60.950 82.890 60.980 ;
        RECT 83.220 60.950 83.880 60.980 ;
        RECT 84.210 60.950 84.870 60.980 ;
        RECT 85.200 60.950 85.860 60.980 ;
        RECT 86.190 60.950 86.850 60.980 ;
        RECT 87.180 60.950 87.840 60.980 ;
        RECT 88.170 60.950 88.830 60.980 ;
        RECT 89.160 60.950 89.820 60.980 ;
        RECT 90.150 60.950 90.810 60.980 ;
        RECT 91.140 60.950 91.800 60.980 ;
        RECT 92.130 60.950 92.790 60.980 ;
        RECT 93.120 60.950 93.780 60.980 ;
        RECT 94.110 60.950 94.770 60.980 ;
        RECT 95.100 60.950 95.760 60.980 ;
        RECT 96.090 60.950 96.750 60.980 ;
        RECT 97.080 60.950 97.740 60.980 ;
        RECT 98.070 60.950 98.730 60.980 ;
        RECT 99.060 60.950 99.720 60.980 ;
        RECT 100.050 60.950 100.710 60.980 ;
        RECT 101.040 60.950 101.700 60.980 ;
        RECT 102.030 60.950 102.690 60.980 ;
        RECT 103.020 60.950 103.680 60.980 ;
        RECT 104.010 60.950 104.670 60.980 ;
        RECT 105.000 60.950 105.660 60.980 ;
        RECT 105.990 60.950 106.650 60.980 ;
        RECT 106.980 60.950 107.640 60.980 ;
        RECT 107.970 60.950 108.630 60.980 ;
        RECT 108.960 60.950 109.620 60.980 ;
        RECT 109.950 60.950 110.610 60.980 ;
        RECT 110.940 60.950 111.600 60.980 ;
        RECT 79.100 60.800 111.600 60.950 ;
        RECT 78.250 58.300 78.650 58.700 ;
        RECT 45.600 40.150 78.100 40.300 ;
        RECT 45.600 40.110 46.260 40.150 ;
        RECT 46.590 40.110 47.250 40.150 ;
        RECT 47.580 40.110 48.240 40.150 ;
        RECT 48.570 40.110 49.230 40.150 ;
        RECT 49.560 40.110 50.220 40.150 ;
        RECT 50.550 40.110 51.210 40.150 ;
        RECT 51.540 40.110 52.200 40.150 ;
        RECT 52.530 40.110 53.190 40.150 ;
        RECT 53.520 40.110 54.180 40.150 ;
        RECT 54.510 40.110 55.170 40.150 ;
        RECT 55.500 40.110 56.160 40.150 ;
        RECT 56.490 40.110 57.150 40.150 ;
        RECT 57.480 40.110 58.140 40.150 ;
        RECT 58.470 40.110 59.130 40.150 ;
        RECT 59.460 40.110 60.120 40.150 ;
        RECT 60.450 40.110 61.110 40.150 ;
        RECT 61.440 40.110 62.100 40.150 ;
        RECT 62.430 40.110 63.090 40.150 ;
        RECT 63.420 40.110 64.080 40.150 ;
        RECT 64.410 40.110 65.070 40.150 ;
        RECT 65.400 40.110 66.060 40.150 ;
        RECT 66.390 40.110 67.050 40.150 ;
        RECT 67.380 40.110 68.040 40.150 ;
        RECT 68.370 40.110 69.030 40.150 ;
        RECT 69.360 40.110 70.020 40.150 ;
        RECT 70.350 40.110 71.010 40.150 ;
        RECT 71.340 40.110 72.000 40.150 ;
        RECT 72.330 40.110 72.990 40.150 ;
        RECT 73.320 40.110 73.980 40.150 ;
        RECT 74.310 40.110 74.970 40.150 ;
        RECT 75.300 40.110 75.960 40.150 ;
        RECT 76.290 40.110 76.950 40.150 ;
        RECT 49.790 39.800 72.760 39.830 ;
        RECT 77.400 39.800 77.800 40.000 ;
        RECT 49.790 39.650 77.800 39.800 ;
        RECT 49.790 39.600 72.760 39.650 ;
        RECT 77.400 39.600 77.800 39.650 ;
        RECT 77.950 39.050 78.100 40.150 ;
        RECT 77.550 38.500 78.100 39.050 ;
        RECT 79.100 40.300 79.250 60.800 ;
        RECT 80.250 60.750 80.910 60.800 ;
        RECT 81.240 60.750 81.900 60.800 ;
        RECT 82.230 60.750 82.890 60.800 ;
        RECT 83.220 60.750 83.880 60.800 ;
        RECT 84.210 60.750 84.870 60.800 ;
        RECT 85.200 60.750 85.860 60.800 ;
        RECT 86.190 60.750 86.850 60.800 ;
        RECT 87.180 60.750 87.840 60.800 ;
        RECT 88.170 60.750 88.830 60.800 ;
        RECT 89.160 60.750 89.820 60.800 ;
        RECT 90.150 60.750 90.810 60.800 ;
        RECT 91.140 60.750 91.800 60.800 ;
        RECT 92.130 60.750 92.790 60.800 ;
        RECT 93.120 60.750 93.780 60.800 ;
        RECT 94.110 60.750 94.770 60.800 ;
        RECT 95.100 60.750 95.760 60.800 ;
        RECT 96.090 60.750 96.750 60.800 ;
        RECT 97.080 60.750 97.740 60.800 ;
        RECT 98.070 60.750 98.730 60.800 ;
        RECT 99.060 60.750 99.720 60.800 ;
        RECT 100.050 60.750 100.710 60.800 ;
        RECT 101.040 60.750 101.700 60.800 ;
        RECT 102.030 60.750 102.690 60.800 ;
        RECT 103.020 60.750 103.680 60.800 ;
        RECT 104.010 60.750 104.670 60.800 ;
        RECT 105.000 60.750 105.660 60.800 ;
        RECT 105.990 60.750 106.650 60.800 ;
        RECT 106.980 60.750 107.640 60.800 ;
        RECT 107.970 60.750 108.630 60.800 ;
        RECT 108.960 60.750 109.620 60.800 ;
        RECT 109.950 60.750 110.610 60.800 ;
        RECT 110.940 60.750 111.600 60.800 ;
        RECT 112.250 59.550 112.400 61.300 ;
        RECT 112.000 59.150 112.400 59.550 ;
        RECT 111.700 58.850 112.750 59.000 ;
        RECT 79.450 58.450 79.850 58.700 ;
        RECT 111.700 58.450 111.850 58.850 ;
        RECT 79.450 58.300 111.850 58.450 ;
        RECT 112.000 58.300 112.400 58.700 ;
        RECT 79.400 42.965 79.630 58.125 ;
        RECT 80.000 57.565 80.150 58.300 ;
        RECT 82.000 57.565 82.150 58.300 ;
        RECT 83.950 57.565 84.100 58.300 ;
        RECT 85.950 57.565 86.100 58.300 ;
        RECT 87.950 57.565 88.100 58.300 ;
        RECT 89.900 57.565 90.050 58.300 ;
        RECT 91.900 57.565 92.050 58.300 ;
        RECT 93.850 57.565 94.000 58.300 ;
        RECT 95.850 57.565 96.000 58.300 ;
        RECT 97.850 57.565 98.000 58.300 ;
        RECT 99.800 57.565 99.950 58.300 ;
        RECT 101.800 57.565 101.950 58.300 ;
        RECT 103.750 57.565 103.900 58.300 ;
        RECT 105.750 57.565 105.900 58.300 ;
        RECT 107.750 57.565 107.900 58.300 ;
        RECT 109.700 57.565 109.850 58.300 ;
        RECT 111.700 57.565 111.850 58.300 ;
        RECT 112.250 58.125 112.400 58.300 ;
        RECT 79.970 43.525 80.200 57.565 ;
        RECT 80.960 43.525 81.190 57.565 ;
        RECT 81.950 43.525 82.180 57.565 ;
        RECT 82.940 43.525 83.170 57.565 ;
        RECT 83.930 43.525 84.160 57.565 ;
        RECT 84.920 43.525 85.150 57.565 ;
        RECT 85.910 43.525 86.140 57.565 ;
        RECT 86.900 43.525 87.130 57.565 ;
        RECT 87.890 43.525 88.120 57.565 ;
        RECT 88.880 43.525 89.110 57.565 ;
        RECT 89.870 43.525 90.100 57.565 ;
        RECT 90.860 43.525 91.090 57.565 ;
        RECT 91.850 43.525 92.080 57.565 ;
        RECT 92.840 43.525 93.070 57.565 ;
        RECT 93.830 43.525 94.060 57.565 ;
        RECT 94.820 43.525 95.050 57.565 ;
        RECT 95.810 43.525 96.040 57.565 ;
        RECT 96.800 43.525 97.030 57.565 ;
        RECT 97.790 43.525 98.020 57.565 ;
        RECT 98.780 43.525 99.010 57.565 ;
        RECT 99.770 43.525 100.000 57.565 ;
        RECT 100.760 43.525 100.990 57.565 ;
        RECT 101.750 43.525 101.980 57.565 ;
        RECT 102.740 43.525 102.970 57.565 ;
        RECT 103.730 43.525 103.960 57.565 ;
        RECT 104.720 43.525 104.950 57.565 ;
        RECT 105.710 43.525 105.940 57.565 ;
        RECT 106.700 43.525 106.930 57.565 ;
        RECT 107.690 43.525 107.920 57.565 ;
        RECT 108.680 43.525 108.910 57.565 ;
        RECT 109.670 43.525 109.900 57.565 ;
        RECT 110.660 43.525 110.890 57.565 ;
        RECT 111.650 43.525 111.880 57.565 ;
        RECT 81.000 42.800 81.150 43.525 ;
        RECT 83.000 42.800 83.150 43.525 ;
        RECT 84.950 42.800 85.100 43.525 ;
        RECT 86.950 42.800 87.100 43.525 ;
        RECT 88.900 42.800 89.050 43.525 ;
        RECT 90.900 42.800 91.050 43.525 ;
        RECT 92.900 42.800 93.050 43.525 ;
        RECT 94.850 42.800 95.000 43.525 ;
        RECT 96.850 42.800 97.000 43.525 ;
        RECT 98.800 42.800 98.950 43.525 ;
        RECT 100.800 42.800 100.950 43.525 ;
        RECT 102.750 42.800 102.900 43.525 ;
        RECT 104.750 42.800 104.900 43.525 ;
        RECT 106.750 42.800 106.900 43.525 ;
        RECT 108.700 42.800 108.850 43.525 ;
        RECT 110.700 42.800 110.850 43.525 ;
        RECT 112.220 42.965 112.450 58.125 ;
        RECT 79.400 42.650 110.850 42.800 ;
        RECT 79.400 42.400 79.800 42.650 ;
        RECT 80.250 40.300 80.910 40.340 ;
        RECT 81.240 40.300 81.900 40.340 ;
        RECT 82.230 40.300 82.890 40.340 ;
        RECT 83.220 40.300 83.880 40.340 ;
        RECT 84.210 40.300 84.870 40.340 ;
        RECT 85.200 40.300 85.860 40.340 ;
        RECT 86.190 40.300 86.850 40.340 ;
        RECT 87.180 40.300 87.840 40.340 ;
        RECT 88.170 40.300 88.830 40.340 ;
        RECT 89.160 40.300 89.820 40.340 ;
        RECT 90.150 40.300 90.810 40.340 ;
        RECT 91.140 40.300 91.800 40.340 ;
        RECT 92.130 40.300 92.790 40.340 ;
        RECT 93.120 40.300 93.780 40.340 ;
        RECT 94.110 40.300 94.770 40.340 ;
        RECT 95.100 40.300 95.760 40.340 ;
        RECT 96.090 40.300 96.750 40.340 ;
        RECT 97.080 40.300 97.740 40.340 ;
        RECT 98.070 40.300 98.730 40.340 ;
        RECT 99.060 40.300 99.720 40.340 ;
        RECT 100.050 40.300 100.710 40.340 ;
        RECT 101.040 40.300 101.700 40.340 ;
        RECT 102.030 40.300 102.690 40.340 ;
        RECT 103.020 40.300 103.680 40.340 ;
        RECT 104.010 40.300 104.670 40.340 ;
        RECT 105.000 40.300 105.660 40.340 ;
        RECT 105.990 40.300 106.650 40.340 ;
        RECT 106.980 40.300 107.640 40.340 ;
        RECT 107.970 40.300 108.630 40.340 ;
        RECT 108.960 40.300 109.620 40.340 ;
        RECT 109.950 40.300 110.610 40.340 ;
        RECT 110.940 40.300 111.600 40.340 ;
        RECT 79.100 40.150 111.600 40.300 ;
        RECT 79.100 39.050 79.250 40.150 ;
        RECT 80.250 40.110 80.910 40.150 ;
        RECT 81.240 40.110 81.900 40.150 ;
        RECT 82.230 40.110 82.890 40.150 ;
        RECT 83.220 40.110 83.880 40.150 ;
        RECT 84.210 40.110 84.870 40.150 ;
        RECT 85.200 40.110 85.860 40.150 ;
        RECT 86.190 40.110 86.850 40.150 ;
        RECT 87.180 40.110 87.840 40.150 ;
        RECT 88.170 40.110 88.830 40.150 ;
        RECT 89.160 40.110 89.820 40.150 ;
        RECT 90.150 40.110 90.810 40.150 ;
        RECT 91.140 40.110 91.800 40.150 ;
        RECT 92.130 40.110 92.790 40.150 ;
        RECT 93.120 40.110 93.780 40.150 ;
        RECT 94.110 40.110 94.770 40.150 ;
        RECT 95.100 40.110 95.760 40.150 ;
        RECT 96.090 40.110 96.750 40.150 ;
        RECT 97.080 40.110 97.740 40.150 ;
        RECT 98.070 40.110 98.730 40.150 ;
        RECT 99.060 40.110 99.720 40.150 ;
        RECT 100.050 40.110 100.710 40.150 ;
        RECT 101.040 40.110 101.700 40.150 ;
        RECT 102.030 40.110 102.690 40.150 ;
        RECT 103.020 40.110 103.680 40.150 ;
        RECT 104.010 40.110 104.670 40.150 ;
        RECT 105.000 40.110 105.660 40.150 ;
        RECT 105.990 40.110 106.650 40.150 ;
        RECT 106.980 40.110 107.640 40.150 ;
        RECT 107.970 40.110 108.630 40.150 ;
        RECT 108.960 40.110 109.620 40.150 ;
        RECT 109.950 40.110 110.610 40.150 ;
        RECT 110.940 40.110 111.600 40.150 ;
        RECT 79.400 39.750 79.800 40.000 ;
        RECT 84.440 39.800 107.410 39.830 ;
        RECT 112.250 39.800 112.400 42.965 ;
        RECT 84.440 39.750 112.400 39.800 ;
        RECT 79.400 39.650 112.400 39.750 ;
        RECT 79.400 39.600 107.410 39.650 ;
        RECT 112.600 39.450 112.750 58.850 ;
        RECT 79.100 38.500 79.650 39.050 ;
        RECT 112.350 38.900 112.900 39.450 ;
        RECT 77.550 37.650 78.100 38.200 ;
        RECT 77.950 2.150 78.100 37.650 ;
        RECT 79.100 37.650 79.650 38.200 ;
        RECT 79.100 2.850 79.250 37.650 ;
        RECT 79.100 2.700 113.700 2.850 ;
        RECT 113.150 2.300 113.700 2.700 ;
        RECT 77.950 2.000 133.050 2.150 ;
        RECT 132.500 1.600 133.050 2.000 ;
      LAYER met2 ;
        RECT 1.000 220.750 3.000 222.750 ;
        RECT 6.000 191.000 8.000 193.000 ;
        RECT 69.750 189.500 70.150 189.750 ;
        RECT 72.800 189.500 73.200 189.750 ;
        RECT 17.550 189.000 17.950 189.400 ;
        RECT 69.750 189.350 73.200 189.500 ;
        RECT 17.550 178.750 17.700 189.000 ;
        RECT 82.550 188.650 82.950 189.050 ;
        RECT 32.200 188.150 32.600 188.400 ;
        RECT 33.350 188.150 33.750 188.400 ;
        RECT 32.200 188.000 59.600 188.150 ;
        RECT 58.850 183.600 59.250 184.000 ;
        RECT 42.050 182.900 42.450 183.300 ;
        RECT 37.500 181.050 37.900 181.300 ;
        RECT 39.350 181.050 39.750 181.450 ;
        RECT 40.300 181.050 40.700 181.300 ;
        RECT 37.500 180.900 40.700 181.050 ;
        RECT 42.050 180.900 42.200 182.900 ;
        RECT 47.950 181.050 48.350 181.300 ;
        RECT 49.800 181.050 50.200 181.450 ;
        RECT 50.750 181.050 51.150 181.300 ;
        RECT 47.950 180.900 51.150 181.050 ;
        RECT 42.050 180.500 42.450 180.900 ;
        RECT 17.550 178.350 17.950 178.750 ;
        RECT 17.550 175.950 17.700 178.350 ;
        RECT 17.550 175.550 17.950 175.950 ;
        RECT 22.050 175.700 22.450 175.850 ;
        RECT 20.600 175.450 22.450 175.700 ;
        RECT 20.600 175.300 21.000 175.450 ;
        RECT 16.600 174.250 19.800 174.400 ;
        RECT 16.600 174.000 17.000 174.250 ;
        RECT 17.850 173.850 18.250 174.250 ;
        RECT 19.400 174.000 19.800 174.250 ;
        RECT 27.050 174.300 27.450 174.550 ;
        RECT 28.900 174.300 29.300 174.700 ;
        RECT 29.850 174.300 30.250 174.550 ;
        RECT 27.050 174.150 30.250 174.300 ;
        RECT 37.500 171.550 37.900 171.800 ;
        RECT 38.450 171.550 38.850 171.950 ;
        RECT 40.300 171.550 40.700 171.800 ;
        RECT 37.500 171.400 40.700 171.550 ;
        RECT 47.950 171.550 48.350 171.800 ;
        RECT 49.050 171.550 49.450 171.950 ;
        RECT 50.750 171.550 51.150 171.800 ;
        RECT 47.950 171.400 51.150 171.550 ;
        RECT 31.050 169.800 31.450 170.050 ;
        RECT 37.500 169.850 37.900 170.100 ;
        RECT 39.350 169.850 39.750 170.250 ;
        RECT 40.300 169.850 40.700 170.100 ;
        RECT 31.050 169.650 32.100 169.800 ;
        RECT 37.500 169.700 40.700 169.850 ;
        RECT 47.950 169.850 48.350 170.100 ;
        RECT 49.800 169.850 50.200 170.250 ;
        RECT 50.750 169.850 51.150 170.100 ;
        RECT 47.950 169.700 51.150 169.850 ;
        RECT 16.600 164.650 17.000 164.900 ;
        RECT 17.550 164.650 17.950 165.050 ;
        RECT 19.400 164.650 19.800 164.900 ;
        RECT 27.050 164.800 27.450 165.050 ;
        RECT 28.000 164.800 28.400 165.200 ;
        RECT 29.850 164.800 30.250 165.050 ;
        RECT 27.050 164.650 30.250 164.800 ;
        RECT 16.600 164.500 19.800 164.650 ;
        RECT 16.600 162.950 17.000 163.200 ;
        RECT 18.100 162.950 18.500 163.350 ;
        RECT 19.400 162.950 19.800 163.200 ;
        RECT 27.050 163.100 27.450 163.350 ;
        RECT 28.900 163.100 29.300 163.500 ;
        RECT 29.850 163.100 30.250 163.350 ;
        RECT 27.050 162.950 30.250 163.100 ;
        RECT 16.600 162.800 19.800 162.950 ;
        RECT 31.950 159.600 32.100 169.650 ;
        RECT 49.200 159.900 49.600 160.150 ;
        RECT 58.850 159.900 59.000 183.600 ;
        RECT 49.200 159.750 59.000 159.900 ;
        RECT 59.450 159.900 59.600 188.000 ;
        RECT 59.750 183.600 60.150 184.000 ;
        RECT 60.400 178.650 60.800 179.050 ;
        RECT 60.650 177.250 60.800 178.650 ;
        RECT 82.800 178.250 82.950 188.650 ;
        RECT 62.550 177.550 62.950 177.950 ;
        RECT 82.550 177.850 82.950 178.250 ;
        RECT 62.550 177.400 70.200 177.550 ;
        RECT 60.650 177.100 69.900 177.250 ;
        RECT 60.350 165.750 60.750 166.150 ;
        RECT 69.750 165.950 69.900 177.100 ;
        RECT 70.050 166.350 70.200 177.400 ;
        RECT 82.800 168.200 82.950 177.850 ;
        RECT 82.800 168.050 113.900 168.200 ;
        RECT 82.800 167.450 82.950 168.050 ;
        RECT 82.550 167.050 82.950 167.450 ;
        RECT 87.100 167.150 87.650 167.700 ;
        RECT 113.750 167.600 113.900 168.050 ;
        RECT 113.750 167.050 114.300 167.600 ;
        RECT 115.400 167.050 115.950 167.600 ;
        RECT 82.800 166.350 82.950 167.050 ;
        RECT 115.400 166.900 115.550 167.050 ;
        RECT 70.050 166.200 82.950 166.350 ;
        RECT 87.950 166.750 115.550 166.900 ;
        RECT 69.750 165.800 84.900 165.950 ;
        RECT 60.350 163.650 60.500 165.750 ;
        RECT 84.750 165.100 84.900 165.800 ;
        RECT 87.950 165.100 88.100 166.750 ;
        RECT 84.500 164.950 88.100 165.100 ;
        RECT 84.500 164.700 84.900 164.950 ;
        RECT 60.350 163.250 60.750 163.650 ;
        RECT 84.750 161.900 84.900 164.700 ;
        RECT 84.500 161.500 84.900 161.900 ;
        RECT 64.500 159.900 64.900 160.150 ;
        RECT 59.450 159.750 64.900 159.900 ;
        RECT 31.950 159.450 51.800 159.600 ;
        RECT 31.600 159.050 32.000 159.300 ;
        RECT 31.600 158.900 51.500 159.050 ;
        RECT 51.350 158.400 51.500 158.900 ;
        RECT 51.650 158.700 51.800 159.450 ;
        RECT 51.950 159.300 62.650 159.450 ;
        RECT 51.950 159.050 52.350 159.300 ;
        RECT 62.250 159.050 62.650 159.300 ;
        RECT 84.750 158.700 84.900 161.500 ;
        RECT 147.000 161.000 149.000 163.000 ;
        RECT 51.650 158.550 52.650 158.700 ;
        RECT 51.350 158.250 51.600 158.400 ;
        RECT 39.900 158.000 40.950 158.150 ;
        RECT 39.900 157.750 40.300 158.000 ;
        RECT 16.600 153.500 17.000 153.750 ;
        RECT 17.550 153.500 17.950 153.900 ;
        RECT 19.400 153.500 19.800 153.750 ;
        RECT 16.600 153.350 19.800 153.500 ;
        RECT 27.050 153.600 27.450 153.850 ;
        RECT 28.000 153.600 28.400 154.000 ;
        RECT 29.850 153.600 30.250 153.850 ;
        RECT 27.050 153.450 30.250 153.600 ;
        RECT 16.600 151.850 17.000 152.100 ;
        RECT 18.100 151.850 18.500 152.250 ;
        RECT 19.400 151.850 19.800 152.100 ;
        RECT 16.600 151.700 19.800 151.850 ;
        RECT 27.050 151.950 27.450 152.200 ;
        RECT 28.900 151.950 29.300 152.350 ;
        RECT 29.850 151.950 30.250 152.200 ;
        RECT 27.050 151.800 30.250 151.950 ;
        RECT 40.800 149.250 40.950 158.000 ;
        RECT 39.850 149.100 40.950 149.250 ;
        RECT 39.850 148.850 40.250 149.100 ;
        RECT 16.600 142.300 17.000 142.550 ;
        RECT 17.550 142.300 17.950 142.700 ;
        RECT 19.400 142.300 19.800 142.550 ;
        RECT 16.600 142.150 19.800 142.300 ;
        RECT 27.050 142.400 27.450 142.650 ;
        RECT 28.000 142.400 28.400 142.800 ;
        RECT 29.850 142.400 30.250 142.650 ;
        RECT 27.050 142.250 30.250 142.400 ;
        RECT 16.600 140.600 17.000 140.850 ;
        RECT 18.100 140.600 18.500 141.000 ;
        RECT 19.400 140.600 19.800 140.850 ;
        RECT 27.050 140.750 27.450 141.000 ;
        RECT 28.900 140.750 29.300 141.150 ;
        RECT 29.850 140.750 30.250 141.000 ;
        RECT 27.050 140.600 30.250 140.750 ;
        RECT 16.600 140.450 19.800 140.600 ;
        RECT 39.900 140.150 40.300 140.400 ;
        RECT 40.800 140.150 40.950 149.100 ;
        RECT 39.900 140.000 40.950 140.150 ;
        RECT 40.800 138.200 40.950 140.000 ;
        RECT 39.900 138.050 40.950 138.200 ;
        RECT 39.900 137.800 40.300 138.050 ;
        RECT 32.000 133.550 32.400 133.950 ;
        RECT 32.000 132.900 32.150 133.550 ;
        RECT 32.000 132.500 32.400 132.900 ;
        RECT 17.550 131.500 17.950 131.900 ;
        RECT 17.550 130.700 17.700 131.500 ;
        RECT 17.550 130.300 17.950 130.700 ;
        RECT 40.800 129.500 40.950 138.050 ;
        RECT 39.900 129.350 40.950 129.500 ;
        RECT 39.900 129.100 40.300 129.350 ;
        RECT 17.550 127.800 17.950 128.200 ;
        RECT 27.600 127.800 28.000 128.050 ;
        RECT 29.450 127.800 29.850 128.050 ;
        RECT 17.550 127.350 17.700 127.800 ;
        RECT 27.600 127.650 29.850 127.800 ;
        RECT 40.800 127.350 40.950 129.350 ;
        RECT 17.550 126.950 17.950 127.350 ;
        RECT 39.900 127.200 40.950 127.350 ;
        RECT 39.900 126.950 40.300 127.200 ;
        RECT 20.550 117.900 20.950 118.100 ;
        RECT 20.550 117.750 23.050 117.900 ;
        RECT 20.550 117.700 20.950 117.750 ;
        RECT 22.650 117.500 23.050 117.750 ;
        RECT 18.220 116.300 18.720 116.600 ;
        RECT 26.920 116.300 27.420 116.600 ;
        RECT 18.220 116.100 27.420 116.300 ;
        RECT 38.020 116.300 38.520 116.600 ;
        RECT 39.550 116.300 39.950 116.500 ;
        RECT 38.020 116.100 40.020 116.300 ;
        RECT 13.320 115.700 40.020 115.900 ;
        RECT 13.320 115.400 13.820 115.700 ;
        RECT 15.820 115.400 16.320 115.700 ;
        RECT 21.720 115.400 22.220 115.700 ;
        RECT 24.120 115.400 24.620 115.700 ;
        RECT 30.120 115.000 30.620 115.700 ;
        RECT 32.520 115.000 33.020 115.700 ;
        RECT 34.920 115.000 35.420 115.700 ;
        RECT 37.320 115.000 37.820 115.700 ;
        RECT 39.520 115.400 40.020 115.700 ;
        RECT 44.120 113.400 49.020 113.600 ;
        RECT 44.120 113.100 44.620 113.400 ;
        RECT 48.820 108.600 49.020 113.400 ;
        RECT 48.520 108.100 49.020 108.600 ;
        RECT 48.520 107.200 49.020 107.700 ;
        RECT 19.720 106.000 20.220 106.300 ;
        RECT 24.620 106.000 25.120 106.300 ;
        RECT 19.720 105.800 25.120 106.000 ;
        RECT 48.820 105.600 49.020 107.200 ;
        RECT 13.320 105.400 49.020 105.600 ;
        RECT 13.320 105.100 13.820 105.400 ;
        RECT 15.720 105.100 16.220 105.400 ;
        RECT 18.120 105.100 18.620 105.400 ;
        RECT 20.620 105.100 21.120 105.400 ;
        RECT 23.020 105.100 23.520 105.400 ;
        RECT 25.520 105.100 26.020 105.400 ;
        RECT 27.920 105.100 28.420 105.400 ;
        RECT 30.320 105.100 30.820 105.400 ;
        RECT 32.720 105.100 33.220 105.400 ;
        RECT 48.620 103.600 49.120 104.100 ;
        RECT 48.920 102.800 49.120 103.600 ;
        RECT 44.220 102.600 49.120 102.800 ;
        RECT 44.220 102.300 44.720 102.600 ;
        RECT 43.520 101.300 44.020 101.800 ;
        RECT 43.820 99.500 44.020 101.300 ;
        RECT 44.520 100.600 44.720 102.300 ;
        RECT 44.220 100.100 44.720 100.600 ;
        RECT 43.520 99.000 44.020 99.500 ;
        RECT 43.820 97.100 44.020 99.000 ;
        RECT 44.520 98.300 44.720 100.100 ;
        RECT 44.220 97.800 44.720 98.300 ;
        RECT 43.520 96.600 44.020 97.100 ;
        RECT 12.320 96.200 12.820 96.500 ;
        RECT 14.820 96.200 15.320 96.500 ;
        RECT 17.220 96.200 17.720 96.500 ;
        RECT 19.620 96.200 20.120 96.500 ;
        RECT 22.020 96.200 22.520 96.500 ;
        RECT 24.520 96.200 25.020 96.500 ;
        RECT 26.920 96.200 27.420 96.500 ;
        RECT 29.420 96.200 29.920 96.500 ;
        RECT 31.820 96.200 32.320 96.500 ;
        RECT 34.120 96.200 34.620 96.500 ;
        RECT 12.320 96.000 34.620 96.200 ;
        RECT 44.400 95.000 44.950 95.550 ;
        RECT 51.450 94.500 51.600 158.250 ;
        RECT 52.500 136.150 52.650 158.550 ;
        RECT 84.500 158.300 84.900 158.700 ;
        RECT 73.300 149.450 73.700 149.850 ;
        RECT 52.500 136.000 59.500 136.150 ;
        RECT 59.350 132.650 59.500 136.000 ;
        RECT 73.300 132.950 73.450 149.450 ;
        RECT 73.600 145.350 83.600 145.500 ;
        RECT 73.600 145.100 74.000 145.350 ;
        RECT 83.200 145.100 83.600 145.350 ;
        RECT 78.550 134.600 78.950 134.850 ;
        RECT 78.250 134.450 78.950 134.600 ;
        RECT 78.250 133.150 78.400 134.450 ;
        RECT 78.550 133.850 78.950 134.250 ;
        RECT 78.800 133.150 78.950 133.850 ;
        RECT 59.900 132.800 73.450 132.950 ;
        RECT 59.350 132.250 59.750 132.650 ;
        RECT 59.900 131.750 60.050 132.800 ;
        RECT 78.000 132.750 78.400 133.150 ;
        RECT 78.550 132.750 78.950 133.150 ;
        RECT 60.200 132.400 60.600 132.650 ;
        RECT 60.200 132.250 97.950 132.400 ;
        RECT 59.650 131.350 60.050 131.750 ;
        RECT 77.350 131.250 77.750 131.500 ;
        RECT 79.450 131.250 79.850 131.500 ;
        RECT 77.350 131.100 79.850 131.250 ;
        RECT 97.800 130.550 97.950 132.250 ;
        RECT 97.800 130.400 108.250 130.550 ;
        RECT 78.550 129.300 78.950 129.550 ;
        RECT 77.600 129.150 78.950 129.300 ;
        RECT 77.600 129.000 77.750 129.150 ;
        RECT 77.350 128.600 77.750 129.000 ;
        RECT 78.250 128.750 78.650 129.000 ;
        RECT 79.450 128.750 79.850 129.000 ;
        RECT 78.250 128.600 79.850 128.750 ;
        RECT 100.550 128.850 100.700 130.400 ;
        RECT 104.150 128.850 104.300 130.400 ;
        RECT 100.550 128.450 100.950 128.850 ;
        RECT 104.150 128.450 104.550 128.850 ;
        RECT 108.100 122.200 108.250 130.400 ;
        RECT 108.100 122.050 109.050 122.200 ;
        RECT 108.650 121.800 109.050 122.050 ;
        RECT 110.750 121.050 111.150 121.300 ;
        RECT 111.650 121.050 112.050 121.300 ;
        RECT 110.750 120.900 112.050 121.050 ;
        RECT 105.650 119.250 106.050 119.650 ;
        RECT 107.400 119.500 107.800 119.900 ;
        RECT 97.850 119.050 98.250 119.150 ;
        RECT 97.850 118.900 99.150 119.050 ;
        RECT 97.850 118.750 98.250 118.900 ;
        RECT 98.750 118.650 99.150 118.900 ;
        RECT 101.450 118.100 101.850 118.300 ;
        RECT 104.150 118.100 104.550 118.300 ;
        RECT 98.100 117.950 104.550 118.100 ;
        RECT 77.400 112.950 77.800 113.200 ;
        RECT 79.400 112.950 79.800 113.200 ;
        RECT 77.400 112.800 79.800 112.950 ;
        RECT 77.350 110.450 77.750 110.700 ;
        RECT 79.450 110.450 79.850 110.700 ;
        RECT 77.350 110.300 79.850 110.450 ;
        RECT 77.350 108.550 79.850 108.700 ;
        RECT 77.350 108.300 77.750 108.550 ;
        RECT 79.450 108.300 79.850 108.550 ;
        RECT 77.350 107.850 77.750 108.100 ;
        RECT 79.450 107.850 79.850 108.100 ;
        RECT 77.350 107.700 79.850 107.850 ;
        RECT 98.100 105.600 98.250 117.950 ;
        RECT 101.450 117.900 101.850 117.950 ;
        RECT 104.150 117.900 104.550 117.950 ;
        RECT 105.650 118.000 105.800 119.250 ;
        RECT 107.650 118.100 107.800 119.500 ;
        RECT 111.650 118.100 111.800 120.900 ;
        RECT 105.650 117.600 106.050 118.000 ;
        RECT 107.650 117.950 111.800 118.100 ;
        RECT 77.350 105.350 77.750 105.600 ;
        RECT 78.250 105.350 78.650 105.600 ;
        RECT 77.350 105.200 78.650 105.350 ;
        RECT 97.500 105.450 98.250 105.600 ;
        RECT 97.500 105.200 97.900 105.450 ;
        RECT 44.400 94.350 51.600 94.500 ;
        RECT 44.400 85.550 44.600 94.350 ;
        RECT 77.400 89.550 77.800 89.800 ;
        RECT 79.400 89.550 79.800 89.800 ;
        RECT 77.400 89.400 79.800 89.550 ;
        RECT 77.350 87.150 79.850 87.300 ;
        RECT 77.350 86.900 77.750 87.150 ;
        RECT 79.450 86.900 79.850 87.150 ;
        RECT 44.200 85.150 44.600 85.550 ;
        RECT 77.400 84.850 79.800 85.000 ;
        RECT 77.400 84.600 77.800 84.850 ;
        RECT 79.400 84.600 79.800 84.850 ;
        RECT 78.550 82.500 78.950 82.750 ;
        RECT 77.600 82.350 78.950 82.500 ;
        RECT 77.600 82.200 77.750 82.350 ;
        RECT 77.350 81.800 77.750 82.200 ;
        RECT 78.250 81.950 78.650 82.200 ;
        RECT 79.450 81.950 79.850 82.200 ;
        RECT 78.250 81.800 79.850 81.950 ;
        RECT 77.400 66.150 79.800 66.300 ;
        RECT 77.400 65.900 77.800 66.150 ;
        RECT 79.400 65.900 79.800 66.150 ;
        RECT 77.700 63.400 78.100 63.800 ;
        RECT 79.100 63.400 79.500 63.800 ;
        RECT 79.100 62.800 79.250 63.400 ;
        RECT 77.400 62.650 79.250 62.800 ;
        RECT 44.750 61.650 45.300 62.200 ;
        RECT 77.400 61.200 77.550 62.650 ;
        RECT 77.700 62.100 78.100 62.500 ;
        RECT 77.950 61.950 78.100 62.100 ;
        RECT 77.950 61.800 79.250 61.950 ;
        RECT 79.100 61.200 79.250 61.800 ;
        RECT 77.400 61.050 78.100 61.200 ;
        RECT 77.700 60.800 78.100 61.050 ;
        RECT 79.100 60.800 79.500 61.200 ;
        RECT 78.550 58.850 78.950 59.250 ;
        RECT 112.000 59.150 112.400 59.550 ;
        RECT 77.350 58.450 77.750 58.700 ;
        RECT 78.250 58.450 78.650 58.700 ;
        RECT 77.350 58.300 78.650 58.450 ;
        RECT 78.800 58.450 78.950 58.850 ;
        RECT 112.250 58.700 112.400 59.150 ;
        RECT 79.450 58.450 79.850 58.700 ;
        RECT 78.800 58.300 79.850 58.450 ;
        RECT 112.000 58.300 112.400 58.700 ;
        RECT 77.400 42.650 79.800 42.800 ;
        RECT 77.400 42.400 77.800 42.650 ;
        RECT 79.400 42.400 79.800 42.650 ;
        RECT 77.400 39.750 77.800 40.000 ;
        RECT 79.400 39.750 79.800 40.000 ;
        RECT 77.400 39.600 79.800 39.750 ;
        RECT 77.550 38.500 78.100 39.050 ;
        RECT 79.100 38.500 79.650 39.050 ;
        RECT 112.350 38.900 112.900 39.450 ;
        RECT 77.550 37.650 78.100 38.200 ;
        RECT 79.100 37.650 79.650 38.200 ;
        RECT 113.150 2.300 113.700 2.850 ;
        RECT 132.500 1.600 133.050 2.150 ;
      LAYER met3 ;
        RECT 1.000 220.750 3.000 222.750 ;
        RECT 6.000 191.000 8.000 193.000 ;
        RECT 87.100 179.800 115.960 190.200 ;
        RECT 87.100 168.200 115.960 178.600 ;
        RECT 87.100 167.150 87.650 167.700 ;
        RECT 113.750 167.050 114.300 167.600 ;
        RECT 115.400 167.050 115.950 167.600 ;
        RECT 147.000 161.000 149.000 163.000 ;
        RECT 44.400 95.000 44.950 95.550 ;
        RECT 12.100 67.300 43.960 94.700 ;
        RECT 113.300 67.300 145.160 94.700 ;
        RECT 12.050 38.700 43.910 66.100 ;
        RECT 44.750 61.650 45.300 62.200 ;
        RECT 12.050 10.100 43.910 37.500 ;
        RECT 45.150 11.600 77.010 39.000 ;
        RECT 77.550 38.500 78.100 39.050 ;
        RECT 79.100 38.500 79.650 39.050 ;
        RECT 77.550 37.650 78.100 38.200 ;
        RECT 79.100 37.650 79.650 38.200 ;
        RECT 80.070 11.580 111.930 38.980 ;
        RECT 112.350 38.900 112.900 39.450 ;
        RECT 113.300 38.700 145.160 66.100 ;
        RECT 113.300 10.100 145.160 37.500 ;
        RECT 113.150 2.300 113.700 2.850 ;
        RECT 132.500 1.600 133.050 2.150 ;
      LAYER met4 ;
        RECT 4.000 224.760 30.670 225.000 ;
        RECT 30.970 224.760 33.430 225.000 ;
        RECT 33.730 224.760 36.190 225.000 ;
        RECT 36.490 224.760 38.950 225.000 ;
        RECT 39.250 224.760 41.710 225.000 ;
        RECT 42.010 224.760 44.470 225.000 ;
        RECT 44.770 224.760 47.230 225.000 ;
        RECT 47.530 224.760 49.990 225.000 ;
        RECT 50.290 224.760 52.750 225.000 ;
        RECT 53.050 224.760 55.510 225.000 ;
        RECT 55.810 224.760 58.270 225.000 ;
        RECT 58.570 224.760 61.030 225.000 ;
        RECT 61.330 224.760 63.790 225.000 ;
        RECT 64.090 224.760 66.550 225.000 ;
        RECT 66.850 224.760 69.310 225.000 ;
        RECT 69.610 224.760 72.070 225.000 ;
        RECT 72.370 224.760 74.830 225.000 ;
        RECT 75.130 224.760 77.590 225.000 ;
        RECT 77.890 224.760 80.350 225.000 ;
        RECT 80.650 224.760 83.110 225.000 ;
        RECT 83.410 224.760 85.870 225.000 ;
        RECT 86.170 224.760 88.630 225.000 ;
        RECT 88.930 224.760 91.390 225.000 ;
        RECT 91.690 224.760 94.150 225.000 ;
        RECT 94.450 224.760 95.000 225.000 ;
        RECT 4.000 224.000 95.000 224.760 ;
        RECT 1.000 220.750 3.000 222.750 ;
        RECT 4.000 220.750 6.000 224.000 ;
        RECT 6.000 191.000 8.000 193.000 ;
        RECT 87.495 180.195 114.105 189.805 ;
        RECT 115.460 180.200 115.940 190.140 ;
        RECT 87.500 178.205 87.800 180.195 ;
        RECT 115.460 179.860 116.550 180.200 ;
        RECT 115.850 179.450 116.550 179.860 ;
        RECT 87.495 168.595 114.105 178.205 ;
        RECT 87.500 167.700 87.800 168.595 ;
        RECT 115.460 168.350 115.940 178.540 ;
        RECT 87.100 167.150 87.800 167.700 ;
        RECT 115.450 167.600 115.950 168.350 ;
        RECT 87.500 132.850 87.800 167.150 ;
        RECT 113.750 167.050 114.300 167.600 ;
        RECT 115.400 167.050 115.950 167.600 ;
        RECT 114.000 166.600 114.300 167.050 ;
        RECT 116.250 166.600 116.550 179.450 ;
        RECT 114.000 166.300 116.550 166.600 ;
        RECT 87.500 132.550 98.400 132.850 ;
        RECT 98.100 131.000 98.400 132.550 ;
        RECT 98.100 130.700 108.700 131.000 ;
        RECT 108.400 123.050 108.700 130.700 ;
        RECT 108.400 122.750 117.100 123.050 ;
        RECT 44.400 95.300 44.950 95.550 ;
        RECT 41.800 95.000 44.950 95.300 ;
        RECT 41.800 94.305 42.100 95.000 ;
        RECT 12.495 67.695 42.105 94.305 ;
        RECT 12.500 65.705 12.800 67.695 ;
        RECT 43.460 67.360 43.940 94.640 ;
        RECT 116.800 94.305 117.100 122.750 ;
        RECT 113.695 67.695 143.305 94.305 ;
        RECT 43.550 66.040 43.850 67.360 ;
        RECT 12.445 39.095 42.055 65.705 ;
        RECT 43.410 61.950 43.890 66.040 ;
        RECT 113.700 65.705 114.000 67.695 ;
        RECT 144.660 67.400 145.140 94.640 ;
        RECT 144.650 65.900 145.150 67.400 ;
        RECT 44.750 61.950 45.300 62.200 ;
        RECT 43.410 61.650 45.300 61.950 ;
        RECT 43.410 39.600 43.890 61.650 ;
        RECT 113.695 40.150 143.305 65.705 ;
        RECT 112.750 40.050 143.305 40.150 ;
        RECT 109.750 39.850 143.305 40.050 ;
        RECT 109.750 39.750 113.050 39.850 ;
        RECT 43.410 39.450 43.950 39.600 ;
        RECT 43.410 39.150 76.950 39.450 ;
        RECT 12.500 37.105 12.800 39.095 ;
        RECT 43.410 38.760 43.900 39.150 ;
        RECT 75.950 38.940 76.950 39.150 ;
        RECT 75.950 38.850 76.990 38.940 ;
        RECT 43.500 37.440 43.900 38.760 ;
        RECT 43.410 37.400 43.900 37.440 ;
        RECT 12.445 10.495 42.055 37.105 ;
        RECT 41.750 9.850 42.050 10.495 ;
        RECT 43.410 10.160 43.890 37.400 ;
        RECT 45.545 12.300 75.155 38.605 ;
        RECT 45.000 11.995 75.155 12.300 ;
        RECT 45.000 9.850 45.850 11.995 ;
        RECT 76.510 11.660 76.990 38.850 ;
        RECT 77.550 38.500 78.100 39.050 ;
        RECT 77.800 38.200 78.100 38.500 ;
        RECT 77.550 37.650 78.100 38.200 ;
        RECT 79.100 38.500 79.650 39.050 ;
        RECT 109.750 38.585 110.750 39.750 ;
        RECT 111.700 38.920 112.900 39.450 ;
        RECT 113.695 39.095 143.305 39.850 ;
        RECT 144.660 39.550 145.140 65.900 ;
        RECT 79.100 38.200 79.400 38.500 ;
        RECT 80.465 38.350 110.750 38.585 ;
        RECT 111.430 38.650 112.900 38.920 ;
        RECT 79.100 37.650 79.650 38.200 ;
        RECT 80.465 12.000 110.075 38.350 ;
        RECT 80.465 11.975 110.750 12.000 ;
        RECT 109.750 11.550 110.750 11.975 ;
        RECT 111.430 11.640 111.910 38.650 ;
        RECT 112.350 38.600 112.900 38.650 ;
        RECT 144.650 38.600 145.150 39.550 ;
        RECT 112.350 38.300 145.150 38.600 ;
        RECT 144.650 37.350 145.150 38.300 ;
        RECT 110.450 11.300 110.750 11.550 ;
        RECT 113.695 11.300 143.305 37.105 ;
        RECT 110.450 11.000 143.305 11.300 ;
        RECT 113.695 10.495 143.305 11.000 ;
        RECT 144.660 10.160 145.140 37.350 ;
        RECT 41.750 9.550 45.850 9.850 ;
        RECT 147.000 3.000 149.000 163.000 ;
        RECT 113.150 2.300 113.700 2.850 ;
        RECT 113.150 1.000 113.650 2.300 ;
        RECT 132.500 1.000 133.050 2.150 ;
        RECT 147.000 1.000 153.000 3.000 ;
        RECT 113.150 0.900 113.170 1.000 ;
  END
END tt_um_rburt16_opamp_3stage
END LIBRARY

