magic
tech sky130A
magscale 1 2
timestamp 1729530615
<< nwell >>
rect -554 -1219 554 1219
<< pmos >>
rect -358 -1000 -158 1000
rect -100 -1000 100 1000
rect 158 -1000 358 1000
<< pdiff >>
rect -416 988 -358 1000
rect -416 -988 -404 988
rect -370 -988 -358 988
rect -416 -1000 -358 -988
rect -158 988 -100 1000
rect -158 -988 -146 988
rect -112 -988 -100 988
rect -158 -1000 -100 -988
rect 100 988 158 1000
rect 100 -988 112 988
rect 146 -988 158 988
rect 100 -1000 158 -988
rect 358 988 416 1000
rect 358 -988 370 988
rect 404 -988 416 988
rect 358 -1000 416 -988
<< pdiffc >>
rect -404 -988 -370 988
rect -146 -988 -112 988
rect 112 -988 146 988
rect 370 -988 404 988
<< nsubdiff >>
rect -518 1149 -422 1183
rect 422 1149 518 1183
rect -518 1087 -484 1149
rect 484 1087 518 1149
rect -518 -1149 -484 -1087
rect 484 -1149 518 -1087
rect -518 -1183 -422 -1149
rect 422 -1183 518 -1149
<< nsubdiffcont >>
rect -422 1149 422 1183
rect -518 -1087 -484 1087
rect 484 -1087 518 1087
rect -422 -1183 422 -1149
<< poly >>
rect -358 1081 -158 1097
rect -358 1047 -342 1081
rect -174 1047 -158 1081
rect -358 1000 -158 1047
rect -100 1081 100 1097
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect -100 1000 100 1047
rect 158 1081 358 1097
rect 158 1047 174 1081
rect 342 1047 358 1081
rect 158 1000 358 1047
rect -358 -1047 -158 -1000
rect -358 -1081 -342 -1047
rect -174 -1081 -158 -1047
rect -358 -1097 -158 -1081
rect -100 -1047 100 -1000
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect -100 -1097 100 -1081
rect 158 -1047 358 -1000
rect 158 -1081 174 -1047
rect 342 -1081 358 -1047
rect 158 -1097 358 -1081
<< polycont >>
rect -342 1047 -174 1081
rect -84 1047 84 1081
rect 174 1047 342 1081
rect -342 -1081 -174 -1047
rect -84 -1081 84 -1047
rect 174 -1081 342 -1047
<< locali >>
rect -518 1149 -422 1183
rect 422 1149 518 1183
rect -518 1087 -484 1149
rect 484 1087 518 1149
rect -358 1047 -342 1081
rect -174 1047 -158 1081
rect -100 1047 -84 1081
rect 84 1047 100 1081
rect 158 1047 174 1081
rect 342 1047 358 1081
rect -404 988 -370 1004
rect -404 -1004 -370 -988
rect -146 988 -112 1004
rect -146 -1004 -112 -988
rect 112 988 146 1004
rect 112 -1004 146 -988
rect 370 988 404 1004
rect 370 -1004 404 -988
rect -358 -1081 -342 -1047
rect -174 -1081 -158 -1047
rect -100 -1081 -84 -1047
rect 84 -1081 100 -1047
rect 158 -1081 174 -1047
rect 342 -1081 358 -1047
rect -518 -1149 -484 -1087
rect 484 -1149 518 -1087
rect -518 -1183 -422 -1149
rect 422 -1183 518 -1149
<< viali >>
rect -342 1047 -174 1081
rect -84 1047 84 1081
rect 174 1047 342 1081
rect -404 -988 -370 988
rect -146 -988 -112 988
rect 112 -988 146 988
rect 370 -988 404 988
rect -342 -1081 -174 -1047
rect -84 -1081 84 -1047
rect 174 -1081 342 -1047
<< metal1 >>
rect -354 1081 -162 1087
rect -354 1047 -342 1081
rect -174 1047 -162 1081
rect -354 1041 -162 1047
rect -96 1081 96 1087
rect -96 1047 -84 1081
rect 84 1047 96 1081
rect -96 1041 96 1047
rect 162 1081 354 1087
rect 162 1047 174 1081
rect 342 1047 354 1081
rect 162 1041 354 1047
rect -410 988 -364 1000
rect -410 -988 -404 988
rect -370 -988 -364 988
rect -410 -1000 -364 -988
rect -152 988 -106 1000
rect -152 -988 -146 988
rect -112 -988 -106 988
rect -152 -1000 -106 -988
rect 106 988 152 1000
rect 106 -988 112 988
rect 146 -988 152 988
rect 106 -1000 152 -988
rect 364 988 410 1000
rect 364 -988 370 988
rect 404 -988 410 988
rect 364 -1000 410 -988
rect -354 -1047 -162 -1041
rect -354 -1081 -342 -1047
rect -174 -1081 -162 -1047
rect -354 -1087 -162 -1081
rect -96 -1047 96 -1041
rect -96 -1081 -84 -1047
rect 84 -1081 96 -1047
rect -96 -1087 96 -1081
rect 162 -1047 354 -1041
rect 162 -1081 174 -1047
rect 342 -1081 354 -1047
rect 162 -1087 354 -1081
<< properties >>
string FIXED_BBOX -501 -1166 501 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
