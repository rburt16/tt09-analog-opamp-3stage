magic
tech sky130A
magscale 1 2
timestamp 1730569394
<< metal1 >>
rect 3200 6600 8520 6640
rect 3200 5840 3240 6600
rect 3300 6120 3340 6600
rect 3400 6400 3500 6420
rect 3400 6340 3420 6400
rect 3480 6340 3500 6400
rect 3400 6240 3500 6340
rect 3680 5840 3720 6600
rect 4380 6540 4480 6560
rect 4380 6480 4400 6540
rect 4460 6480 4480 6540
rect 4380 6460 4480 6480
rect 3900 6400 4000 6420
rect 3900 6340 3920 6400
rect 3980 6340 4000 6400
rect 3900 6240 4000 6340
rect 4380 6280 4420 6460
rect 4380 6240 4520 6280
rect 4380 6140 4420 6240
rect 4280 5840 4320 5880
rect 4860 5840 4900 6600
rect 4980 6120 5020 6600
rect 5080 6400 5180 6420
rect 5080 6340 5100 6400
rect 5160 6340 5180 6400
rect 5080 6240 5180 6340
rect 5360 5840 5400 6600
rect 6120 6540 6220 6560
rect 6120 6480 6140 6540
rect 6200 6480 6220 6540
rect 6120 6460 6220 6480
rect 5560 6400 5660 6420
rect 5560 6340 5580 6400
rect 5640 6340 5660 6400
rect 5560 6280 5660 6340
rect 5560 6240 6100 6280
rect 6160 6240 6220 6460
rect 6060 6140 6100 6240
rect 5960 5840 5980 5880
rect 6540 5840 6580 6600
rect 6660 6120 6700 6600
rect 6760 6400 6860 6420
rect 6760 6340 6780 6400
rect 6840 6340 6860 6400
rect 6760 6240 6860 6340
rect 7020 5840 7060 6600
rect 7240 6400 7340 6420
rect 7240 6340 7260 6400
rect 7320 6340 7340 6400
rect 7240 6240 7340 6340
rect 7500 5840 7540 6600
rect 7620 6120 7660 6600
rect 7720 6400 7820 6420
rect 7720 6340 7740 6400
rect 7800 6340 7820 6400
rect 7720 6240 7820 6340
rect 7980 5840 8020 6600
rect 8340 6540 8440 6560
rect 8340 6480 8360 6540
rect 8420 6480 8440 6540
rect 8340 6460 8440 6480
rect 8200 6400 8300 6420
rect 8200 6340 8220 6400
rect 8280 6340 8300 6400
rect 8200 6240 8300 6340
rect 8380 6140 8420 6460
rect 8480 5260 8520 6600
rect 8640 6400 8740 6420
rect 8640 6340 8660 6400
rect 8720 6340 8740 6400
rect 8640 6320 8740 6340
rect 8580 5540 8620 5700
rect 8700 5680 8740 6320
rect 9560 5940 9660 5960
rect 9560 5880 9580 5940
rect 9640 5880 9660 5940
rect 9560 5860 9660 5880
rect 9560 5780 9600 5860
rect 10360 5540 10400 5700
rect 8580 5500 10700 5540
rect 9800 5320 10620 5360
rect 8480 5220 8640 5260
rect 10260 5200 10540 5240
rect 10500 4960 10540 5200
rect 10440 4940 10540 4960
rect 10440 4900 10460 4940
rect 10240 4880 10460 4900
rect 10520 4880 10540 4940
rect 10240 4860 10540 4880
rect 10580 4780 10620 5320
rect 10340 4760 10620 4780
rect 10340 4740 10460 4760
rect 3580 4600 3820 4640
rect 4060 4600 4420 4640
rect 4660 4580 4700 4640
rect 5260 4600 5500 4640
rect 5740 4600 6100 4640
rect 4660 4540 4860 4580
rect 4680 4480 4780 4500
rect 4680 4440 4700 4480
rect 3280 4420 4700 4440
rect 4760 4420 4780 4480
rect 4820 4480 4860 4540
rect 5660 4480 5760 4500
rect 4820 4440 5280 4480
rect 3280 4400 4780 4420
rect 3280 4120 3320 4400
rect 3400 4340 3500 4360
rect 3400 4280 3420 4340
rect 3480 4280 3500 4340
rect 3400 4220 3500 4280
rect 3780 4120 3820 4400
rect 3880 4340 3980 4360
rect 3880 4280 3900 4340
rect 3960 4280 3980 4340
rect 3880 4220 3980 4280
rect 4260 4120 4300 4400
rect 4360 4340 4460 4360
rect 4360 4280 4380 4340
rect 4440 4280 4460 4340
rect 4360 4220 4460 4280
rect 4740 4120 4780 4400
rect 5240 4360 5280 4440
rect 5660 4420 5680 4480
rect 5740 4440 5760 4480
rect 6340 4440 6380 4640
rect 6940 4620 7180 4660
rect 7420 4440 7460 4640
rect 7900 4600 8140 4640
rect 8600 4520 8640 4720
rect 10440 4700 10460 4740
rect 10520 4740 10620 4760
rect 10520 4700 10540 4740
rect 10440 4680 10540 4700
rect 8720 4520 8760 4620
rect 10660 4520 10700 5500
rect 8600 4480 10700 4520
rect 5740 4420 7220 4440
rect 5660 4400 7220 4420
rect 7420 4400 10400 4440
rect 4860 4340 4960 4360
rect 4860 4280 4880 4340
rect 4940 4280 4960 4340
rect 4860 4220 4960 4280
rect 5240 4340 5440 4360
rect 5240 4320 5360 4340
rect 5240 4120 5280 4320
rect 5340 4280 5360 4320
rect 5420 4280 5440 4340
rect 5340 4220 5440 4280
rect 5720 4120 5760 4400
rect 5840 4340 5940 4360
rect 5840 4280 5860 4340
rect 5920 4280 5940 4340
rect 5840 4220 5940 4280
rect 6200 4120 6240 4400
rect 6320 4340 6420 4360
rect 6320 4280 6340 4340
rect 6400 4280 6420 4340
rect 6320 4220 6420 4280
rect 6700 4120 6740 4400
rect 6800 4340 6900 4360
rect 6800 4280 6820 4340
rect 6880 4280 6900 4340
rect 6800 4220 6900 4280
rect 7180 4120 7220 4400
rect 7280 4340 7380 4360
rect 7280 4280 7300 4340
rect 7360 4280 7380 4340
rect 7280 4220 7380 4280
rect 10360 4220 10400 4400
rect 9640 4180 10400 4220
rect 10360 4080 10400 4180
rect 10460 4040 10560 4060
rect 10460 4000 10480 4040
rect 7680 3620 7720 4000
rect 10380 3980 10480 4000
rect 10540 3980 10560 4040
rect 10380 3960 10560 3980
rect 9580 3780 9680 3800
rect 9580 3760 9600 3780
rect 8880 3720 9600 3760
rect 9660 3720 9680 3780
rect 9580 3700 9680 3720
rect 9720 3720 9760 3860
rect 10600 3720 10640 4480
rect 9720 3680 10640 3720
rect 9440 3580 9540 3600
rect 9440 3560 9460 3580
rect 9360 3520 9460 3560
rect 9520 3520 9540 3580
rect 9360 3500 9540 3520
rect 9720 3460 9760 3680
rect 9440 3420 9760 3460
rect 7560 3360 8120 3400
rect 8960 3380 9480 3420
rect 7560 2940 7600 3360
rect 9580 3340 9680 3360
rect 9580 3300 9600 3340
rect 8880 3280 9600 3300
rect 9660 3280 9680 3340
rect 8880 3260 9680 3280
rect 9440 3120 9540 3140
rect 9440 3100 9460 3120
rect 7680 2940 7720 3100
rect 9360 3060 9460 3100
rect 9520 3060 9540 3120
rect 9360 3040 9540 3060
rect 7560 2900 8120 2940
rect 3200 2520 3300 2540
rect 3200 2460 3220 2520
rect 3280 2480 3300 2520
rect 3280 2460 3400 2480
rect 3200 2440 3400 2460
rect 3580 2400 3620 2620
rect 3700 2520 3800 2540
rect 3700 2460 3720 2520
rect 3780 2480 3800 2520
rect 3780 2460 3900 2480
rect 3700 2440 3900 2460
rect 4060 2400 4100 2620
rect 4180 2520 4280 2540
rect 4180 2460 4200 2520
rect 4260 2480 4280 2520
rect 4260 2460 4380 2480
rect 4180 2440 4380 2460
rect 4540 2400 4580 2620
rect 4660 2520 4760 2540
rect 4660 2460 4680 2520
rect 4740 2480 4760 2520
rect 4740 2460 4880 2480
rect 4660 2440 4880 2460
rect 5040 2400 5080 2620
rect 5140 2520 5240 2540
rect 5140 2460 5160 2520
rect 5220 2480 5240 2520
rect 5520 2480 5560 2620
rect 5220 2460 5560 2480
rect 5140 2440 5560 2460
rect 5640 2520 5740 2540
rect 5640 2460 5660 2520
rect 5720 2480 5740 2520
rect 5720 2460 5840 2480
rect 5640 2440 5840 2460
rect 6000 2400 6040 2620
rect 6120 2520 6220 2540
rect 6120 2460 6140 2520
rect 6200 2480 6220 2520
rect 6200 2460 6320 2480
rect 6120 2440 6320 2460
rect 6480 2400 6520 2620
rect 6620 2520 6720 2540
rect 6620 2460 6640 2520
rect 6700 2480 6720 2520
rect 6700 2460 6820 2480
rect 6620 2440 6820 2460
rect 6980 2400 7020 2620
rect 7100 2520 7200 2540
rect 7100 2460 7120 2520
rect 7180 2480 7200 2520
rect 7180 2460 7320 2480
rect 7100 2440 7320 2460
rect 7460 2400 7500 2620
rect 7560 2540 7600 2900
rect 9580 2880 9680 2900
rect 9580 2840 9600 2880
rect 8880 2820 9600 2840
rect 9660 2820 9680 2880
rect 8880 2800 9680 2820
rect 9440 2640 9540 2660
rect 7680 2540 7720 2640
rect 9440 2620 9460 2640
rect 7560 2520 7720 2540
rect 7560 2460 7580 2520
rect 7640 2480 7720 2520
rect 9360 2580 9460 2620
rect 9520 2580 9540 2640
rect 9360 2560 9540 2580
rect 7640 2460 8120 2480
rect 7560 2440 8120 2460
rect 9360 2400 9400 2560
rect 3580 2360 9400 2400
<< via1 >>
rect 3420 6340 3480 6400
rect 4400 6480 4460 6540
rect 3920 6340 3980 6400
rect 5100 6340 5160 6400
rect 6140 6480 6200 6540
rect 5580 6340 5640 6400
rect 6780 6340 6840 6400
rect 7260 6340 7320 6400
rect 7740 6340 7800 6400
rect 8360 6480 8420 6540
rect 8220 6340 8280 6400
rect 8660 6340 8720 6400
rect 9580 5880 9640 5940
rect 10460 4880 10520 4940
rect 4700 4420 4760 4480
rect 3420 4280 3480 4340
rect 3900 4280 3960 4340
rect 4380 4280 4440 4340
rect 5680 4420 5740 4480
rect 10460 4700 10520 4760
rect 4880 4280 4940 4340
rect 5360 4280 5420 4340
rect 5860 4280 5920 4340
rect 6340 4280 6400 4340
rect 6820 4280 6880 4340
rect 7300 4280 7360 4340
rect 10480 3980 10540 4040
rect 9600 3720 9660 3780
rect 9460 3520 9520 3580
rect 9600 3280 9660 3340
rect 9460 3060 9520 3120
rect 3220 2460 3280 2520
rect 3720 2460 3780 2520
rect 4200 2460 4260 2520
rect 4680 2460 4740 2520
rect 5160 2460 5220 2520
rect 5660 2460 5720 2520
rect 6140 2460 6200 2520
rect 6640 2460 6700 2520
rect 7120 2460 7180 2520
rect 9600 2820 9660 2880
rect 7580 2460 7640 2520
rect 9460 2580 9520 2640
<< metal2 >>
rect 4380 6540 4480 6560
rect 4380 6480 4400 6540
rect 4460 6500 4480 6540
rect 6120 6540 6220 6560
rect 6120 6500 6140 6540
rect 4460 6480 6140 6500
rect 6200 6480 6220 6540
rect 4380 6460 6220 6480
rect 8340 6540 8440 6560
rect 8340 6480 8360 6540
rect 8420 6500 8440 6540
rect 8420 6480 8740 6500
rect 8340 6460 8740 6480
rect 3400 6400 8740 6420
rect 3400 6340 3420 6400
rect 3480 6380 3920 6400
rect 3480 6340 3500 6380
rect 3400 6320 3500 6340
rect 3900 6340 3920 6380
rect 3980 6380 5100 6400
rect 3980 6340 4000 6380
rect 3900 6320 4000 6340
rect 5080 6340 5100 6380
rect 5160 6380 5580 6400
rect 5160 6340 5180 6380
rect 5080 6320 5180 6340
rect 5560 6340 5580 6380
rect 5640 6380 6780 6400
rect 5640 6340 5660 6380
rect 5560 6320 5660 6340
rect 6760 6340 6780 6380
rect 6840 6380 7260 6400
rect 6840 6340 6860 6380
rect 6760 6240 6860 6340
rect 7240 6340 7260 6380
rect 7320 6380 7740 6400
rect 7320 6340 7340 6380
rect 7240 6240 7340 6340
rect 7720 6340 7740 6380
rect 7800 6380 8220 6400
rect 7800 6340 7820 6380
rect 7720 6240 7820 6340
rect 8200 6340 8220 6380
rect 8280 6380 8660 6400
rect 8280 6340 8300 6380
rect 8200 6240 8300 6340
rect 8640 6340 8660 6380
rect 8720 6340 8740 6400
rect 8640 6320 8740 6340
rect 9560 5940 10540 5960
rect 9560 5880 9580 5940
rect 9640 5920 10540 5940
rect 9640 5880 9660 5920
rect 9560 5860 9660 5880
rect 10500 4960 10540 5920
rect 10440 4940 10540 4960
rect 10440 4880 10460 4940
rect 10520 4880 10540 4940
rect 10440 4860 10540 4880
rect 10440 4760 10540 4780
rect 10440 4700 10460 4760
rect 10520 4700 10540 4760
rect 10440 4680 10540 4700
rect 4680 4480 4780 4500
rect 4680 4420 4700 4480
rect 4760 4440 4780 4480
rect 5660 4480 5760 4500
rect 5660 4440 5680 4480
rect 4760 4420 5680 4440
rect 5740 4420 5760 4480
rect 4680 4400 5760 4420
rect 10500 4360 10540 4680
rect 3400 4340 10540 4360
rect 3400 4280 3420 4340
rect 3480 4320 3900 4340
rect 3480 4280 3500 4320
rect 3400 4260 3500 4280
rect 3880 4280 3900 4320
rect 3960 4320 4380 4340
rect 3960 4280 3980 4320
rect 3880 4260 3980 4280
rect 4360 4280 4380 4320
rect 4440 4320 4880 4340
rect 4440 4280 4460 4320
rect 4360 4260 4460 4280
rect 4860 4280 4880 4320
rect 4940 4320 5360 4340
rect 4940 4280 4960 4320
rect 4860 4260 4960 4280
rect 5340 4280 5360 4320
rect 5420 4320 5860 4340
rect 5420 4280 5440 4320
rect 5340 4260 5440 4280
rect 5840 4280 5860 4320
rect 5920 4320 6340 4340
rect 5920 4280 5940 4320
rect 5840 4260 5940 4280
rect 6320 4280 6340 4320
rect 6400 4320 6820 4340
rect 6400 4280 6420 4320
rect 6320 4260 6420 4280
rect 6800 4280 6820 4320
rect 6880 4320 7300 4340
rect 6880 4280 6900 4320
rect 6800 4260 6900 4280
rect 7280 4280 7300 4320
rect 7360 4320 10540 4340
rect 7360 4280 7380 4320
rect 7280 4260 7380 4280
rect 10460 4040 10560 4060
rect 10460 3980 10480 4040
rect 10540 3980 10560 4040
rect 10460 3960 10560 3980
rect 10520 3800 10560 3960
rect 9580 3780 10560 3800
rect 9580 3720 9600 3780
rect 9660 3760 10560 3780
rect 9660 3720 9680 3760
rect 9580 3700 9680 3720
rect 9440 3580 9540 3600
rect 9440 3520 9460 3580
rect 9520 3520 9540 3580
rect 9440 3500 9540 3520
rect 9500 3140 9540 3500
rect 9640 3360 9680 3700
rect 9580 3340 9680 3360
rect 9580 3280 9600 3340
rect 9660 3280 9680 3340
rect 9580 3260 9680 3280
rect 9440 3120 9540 3140
rect 9440 3060 9460 3120
rect 9520 3060 9540 3120
rect 9440 3040 9540 3060
rect 9500 2660 9540 3040
rect 9640 2900 9680 3260
rect 9580 2880 9680 2900
rect 9580 2820 9600 2880
rect 9660 2820 9680 2880
rect 9580 2800 9680 2820
rect 9440 2640 9540 2660
rect 9440 2580 9460 2640
rect 9520 2580 9540 2640
rect 9440 2560 9540 2580
rect 3200 2520 3300 2540
rect 3200 2460 3220 2520
rect 3280 2480 3300 2520
rect 3700 2520 3800 2540
rect 3700 2480 3720 2520
rect 3280 2460 3720 2480
rect 3780 2480 3800 2520
rect 4180 2520 4280 2540
rect 4180 2480 4200 2520
rect 3780 2460 4200 2480
rect 4260 2480 4280 2520
rect 4660 2520 4760 2540
rect 4660 2480 4680 2520
rect 4260 2460 4680 2480
rect 4740 2480 4760 2520
rect 5140 2520 5240 2540
rect 5140 2480 5160 2520
rect 4740 2460 5160 2480
rect 5220 2480 5240 2520
rect 5640 2520 5740 2540
rect 5640 2480 5660 2520
rect 5220 2460 5660 2480
rect 5720 2480 5740 2520
rect 6120 2520 6220 2540
rect 6120 2480 6140 2520
rect 5720 2460 6140 2480
rect 6200 2480 6220 2520
rect 6620 2520 6720 2540
rect 6620 2480 6640 2520
rect 6200 2460 6640 2480
rect 6700 2480 6720 2520
rect 7100 2520 7200 2540
rect 7100 2480 7120 2520
rect 6700 2460 7120 2480
rect 7180 2480 7200 2520
rect 7560 2520 7660 2540
rect 7560 2480 7580 2520
rect 7180 2460 7580 2480
rect 7640 2460 7660 2520
rect 3200 2440 7660 2460
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_0
timestamp 1730569394
transform 1 0 3452 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_1
timestamp 1730569394
transform 1 0 5396 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_2
timestamp 1730569394
transform 1 0 4910 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_3
timestamp 1730569394
transform 1 0 4424 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_4
timestamp 1730569394
transform 1 0 3938 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_5
timestamp 1730569394
transform 1 0 6368 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_6
timestamp 1730569394
transform 1 0 5882 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_7
timestamp 1730569394
transform 1 0 7340 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_92UKLN  sky130_fd_pr__nfet_01v8_92UKLN_8
timestamp 1730569394
transform 1 0 6854 0 1 3399
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_EE6UX6  sky130_fd_pr__nfet_01v8_EE6UX6_0
timestamp 1730569394
transform 1 0 8536 0 1 2699
box -996 -279 996 279
use sky130_fd_pr__nfet_01v8_EE6UX6  sky130_fd_pr__nfet_01v8_EE6UX6_1
timestamp 1730569394
transform 1 0 8536 0 1 3159
box -996 -279 996 279
use sky130_fd_pr__nfet_01v8_QGAK58  sky130_fd_pr__nfet_01v8_QGAK58_0
timestamp 1730569394
transform 0 1 9539 -1 0 4736
box -296 -979 296 979
use sky130_fd_pr__pfet_01v8_L7EPZQ  sky130_fd_pr__pfet_01v8_L7EPZQ_0
timestamp 1730569394
transform 1 0 7776 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_lvt_LBMMZQ  sky130_fd_pr__pfet_01v8_lvt_LBMMZQ_0
timestamp 1730569394
transform 1 0 8255 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_BMAEVH  XM3
timestamp 1730569394
transform 1 0 3456 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_L7EPZQ  XM4
timestamp 1730569394
transform 1 0 5136 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_L7EPZQ  XM6
timestamp 1730569394
transform 1 0 6816 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__nfet_01v8_798YF4  XM7
timestamp 1730569394
transform 1 0 9046 0 1 4079
box -1506 -279 1506 279
use sky130_fd_pr__nfet_01v8_EE6UX6  XM8
timestamp 1730569394
transform 1 0 8536 0 1 3619
box -996 -279 996 279
use sky130_fd_pr__nfet_01v8_lvt_XLZA2Q  XM9
timestamp 1730569394
transform 1 0 4536 0 1 5419
box -296 -979 296 979
use sky130_fd_pr__nfet_01v8_lvt_X6KF3T  XM10
timestamp 1730569394
transform 1 0 6218 0 1 5422
box -296 -979 296 979
use sky130_fd_pr__pfet_01v8_lvt_LHEPZQ  XM11
timestamp 1730569394
transform 1 0 3942 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_lvt_LBMMZQ  XM12
timestamp 1730569394
transform 1 0 5622 0 1 5425
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_lvt_LBMMZQ  XM13
timestamp 1730569394
transform 1 0 7296 0 1 5424
box -296 -984 296 984
use sky130_fd_pr__pfet_01v8_GQTHCS  XM16
timestamp 1730569394
transform 1 0 9456 0 1 5266
box -996 -226 996 226
use sky130_fd_pr__nfet_01v8_N4YVNS  XM18
timestamp 1730569394
transform 1 0 9556 0 1 5721
box -996 -221 996 221
<< end >>
