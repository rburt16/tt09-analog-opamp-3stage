magic
tech sky130A
magscale 1 2
timestamp 1730482424
<< error_p >>
rect -31 4435 31 4441
rect -31 4401 -19 4435
rect -31 4395 31 4401
rect -31 2307 31 2313
rect -31 2273 -19 2307
rect -31 2267 31 2273
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect -31 2159 31 2165
rect -31 71 31 77
rect -31 37 -19 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect -31 -77 31 -71
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect -31 -2205 31 -2199
rect -31 -2273 31 -2267
rect -31 -2307 -19 -2273
rect -31 -2313 31 -2307
rect -31 -4401 31 -4395
rect -31 -4435 -19 -4401
rect -31 -4441 31 -4435
<< nwell >>
rect -231 -4573 231 4573
<< pmoslvt >>
rect -35 2354 35 4354
rect -35 118 35 2118
rect -35 -2118 35 -118
rect -35 -4354 35 -2354
<< pdiff >>
rect -93 4046 -35 4354
rect -93 2662 -81 4046
rect -47 2662 -35 4046
rect -93 2354 -35 2662
rect 35 4046 93 4354
rect 35 2662 47 4046
rect 81 2662 93 4046
rect 35 2354 93 2662
rect -93 1810 -35 2118
rect -93 426 -81 1810
rect -47 426 -35 1810
rect -93 118 -35 426
rect 35 1810 93 2118
rect 35 426 47 1810
rect 81 426 93 1810
rect 35 118 93 426
rect -93 -426 -35 -118
rect -93 -1810 -81 -426
rect -47 -1810 -35 -426
rect -93 -2118 -35 -1810
rect 35 -426 93 -118
rect 35 -1810 47 -426
rect 81 -1810 93 -426
rect 35 -2118 93 -1810
rect -93 -2662 -35 -2354
rect -93 -4046 -81 -2662
rect -47 -4046 -35 -2662
rect -93 -4354 -35 -4046
rect 35 -2662 93 -2354
rect 35 -4046 47 -2662
rect 81 -4046 93 -2662
rect 35 -4354 93 -4046
<< pdiffc >>
rect -81 2662 -47 4046
rect 47 2662 81 4046
rect -81 426 -47 1810
rect 47 426 81 1810
rect -81 -1810 -47 -426
rect 47 -1810 81 -426
rect -81 -4046 -47 -2662
rect 47 -4046 81 -2662
<< nsubdiff >>
rect -195 4503 -69 4537
rect 69 4503 195 4537
rect -195 3109 -161 4503
rect 161 3109 195 4503
rect -195 -4503 -161 -3109
rect 161 -4503 195 -3109
rect -195 -4537 -69 -4503
rect 69 -4537 195 -4503
<< nsubdiffcont >>
rect -69 4503 69 4537
rect -195 -3109 -161 3109
rect 161 -3109 195 3109
rect -69 -4537 69 -4503
<< poly >>
rect -33 4435 33 4451
rect -33 4418 -17 4435
rect -35 4401 -17 4418
rect 17 4418 33 4435
rect 17 4401 35 4418
rect -35 4354 35 4401
rect -35 2307 35 2354
rect -35 2290 -17 2307
rect -33 2273 -17 2290
rect 17 2290 35 2307
rect 17 2273 33 2290
rect -33 2257 33 2273
rect -33 2199 33 2215
rect -33 2182 -17 2199
rect -35 2165 -17 2182
rect 17 2182 33 2199
rect 17 2165 35 2182
rect -35 2118 35 2165
rect -35 71 35 118
rect -35 54 -17 71
rect -33 37 -17 54
rect 17 54 35 71
rect 17 37 33 54
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -54 -17 -37
rect -35 -71 -17 -54
rect 17 -54 33 -37
rect 17 -71 35 -54
rect -35 -118 35 -71
rect -35 -2165 35 -2118
rect -35 -2182 -17 -2165
rect -33 -2199 -17 -2182
rect 17 -2182 35 -2165
rect 17 -2199 33 -2182
rect -33 -2215 33 -2199
rect -33 -2273 33 -2257
rect -33 -2290 -17 -2273
rect -35 -2307 -17 -2290
rect 17 -2290 33 -2273
rect 17 -2307 35 -2290
rect -35 -2354 35 -2307
rect -35 -4401 35 -4354
rect -35 -4418 -17 -4401
rect -33 -4435 -17 -4418
rect 17 -4418 35 -4401
rect 17 -4435 33 -4418
rect -33 -4451 33 -4435
<< polycont >>
rect -17 4401 17 4435
rect -17 2273 17 2307
rect -17 2165 17 2199
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -2199 17 -2165
rect -17 -2307 17 -2273
rect -17 -4435 17 -4401
<< locali >>
rect -195 4503 -113 4537
rect 113 4503 195 4537
rect -195 3152 -161 4503
rect -33 4401 -19 4435
rect 19 4401 33 4435
rect -81 4046 -47 4062
rect -81 2646 -47 2662
rect 47 4046 81 4062
rect 47 2646 81 2662
rect 161 3152 195 4503
rect -33 2273 -19 2307
rect 19 2273 33 2307
rect -33 2165 -19 2199
rect 19 2165 33 2199
rect -81 1810 -47 1826
rect -81 410 -47 426
rect 47 1810 81 1826
rect 47 410 81 426
rect -33 37 -19 71
rect 19 37 33 71
rect -33 -71 -19 -37
rect 19 -71 33 -37
rect -81 -426 -47 -410
rect -81 -1826 -47 -1810
rect 47 -426 81 -410
rect 47 -1826 81 -1810
rect -33 -2199 -19 -2165
rect 19 -2199 33 -2165
rect -33 -2307 -19 -2273
rect 19 -2307 33 -2273
rect -195 -4503 -161 -3152
rect -81 -2662 -47 -2646
rect -81 -4062 -47 -4046
rect 47 -2662 81 -2646
rect 47 -4062 81 -4046
rect -33 -4435 -19 -4401
rect 19 -4435 33 -4401
rect 161 -4503 195 -3152
rect -195 -4537 -113 -4503
rect 113 -4537 195 -4503
<< viali >>
rect -113 4503 -69 4537
rect -69 4503 69 4537
rect 69 4503 113 4537
rect -19 4401 -17 4435
rect -17 4401 17 4435
rect 17 4401 19 4435
rect -195 3109 -161 3152
rect -195 -3109 -161 3109
rect -81 2662 -47 4046
rect 47 2662 81 4046
rect 161 3109 195 3152
rect -19 2273 -17 2307
rect -17 2273 17 2307
rect 17 2273 19 2307
rect -19 2165 -17 2199
rect -17 2165 17 2199
rect 17 2165 19 2199
rect -81 426 -47 1810
rect 47 426 81 1810
rect -19 37 -17 71
rect -17 37 17 71
rect 17 37 19 71
rect -19 -71 -17 -37
rect -17 -71 17 -37
rect 17 -71 19 -37
rect -81 -1810 -47 -426
rect 47 -1810 81 -426
rect -19 -2199 -17 -2165
rect -17 -2199 17 -2165
rect 17 -2199 19 -2165
rect -19 -2307 -17 -2273
rect -17 -2307 17 -2273
rect 17 -2307 19 -2273
rect -195 -3152 -161 -3109
rect -81 -4046 -47 -2662
rect 47 -4046 81 -2662
rect 161 -3109 195 3109
rect 161 -3152 195 -3109
rect -19 -4435 -17 -4401
rect -17 -4435 17 -4401
rect 17 -4435 19 -4401
rect -113 -4537 -69 -4503
rect -69 -4537 69 -4503
rect 69 -4537 113 -4503
<< metal1 >>
rect -125 4537 125 4543
rect -125 4503 -113 4537
rect 113 4503 125 4537
rect -125 4497 125 4503
rect -31 4435 31 4441
rect -31 4401 -19 4435
rect 19 4401 31 4435
rect -31 4395 31 4401
rect -87 4046 -41 4058
rect -201 3152 -155 3164
rect -201 -3152 -195 3152
rect -161 -3152 -155 3152
rect -87 2662 -81 4046
rect -47 2662 -41 4046
rect -87 2650 -41 2662
rect 41 4046 87 4058
rect 41 2662 47 4046
rect 81 2662 87 4046
rect 41 2650 87 2662
rect 155 3152 201 3164
rect -31 2307 31 2313
rect -31 2273 -19 2307
rect 19 2273 31 2307
rect -31 2267 31 2273
rect -31 2199 31 2205
rect -31 2165 -19 2199
rect 19 2165 31 2199
rect -31 2159 31 2165
rect -87 1810 -41 1822
rect -87 426 -81 1810
rect -47 426 -41 1810
rect -87 414 -41 426
rect 41 1810 87 1822
rect 41 426 47 1810
rect 81 426 87 1810
rect 41 414 87 426
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect -87 -426 -41 -414
rect -87 -1810 -81 -426
rect -47 -1810 -41 -426
rect -87 -1822 -41 -1810
rect 41 -426 87 -414
rect 41 -1810 47 -426
rect 81 -1810 87 -426
rect 41 -1822 87 -1810
rect -31 -2165 31 -2159
rect -31 -2199 -19 -2165
rect 19 -2199 31 -2165
rect -31 -2205 31 -2199
rect -31 -2273 31 -2267
rect -31 -2307 -19 -2273
rect 19 -2307 31 -2273
rect -31 -2313 31 -2307
rect -201 -3164 -155 -3152
rect -87 -2662 -41 -2650
rect -87 -4046 -81 -2662
rect -47 -4046 -41 -2662
rect -87 -4058 -41 -4046
rect 41 -2662 87 -2650
rect 41 -4046 47 -2662
rect 81 -4046 87 -2662
rect 155 -3152 161 3152
rect 195 -3152 201 3152
rect 155 -3164 201 -3152
rect 41 -4058 87 -4046
rect -31 -4401 31 -4395
rect -31 -4435 -19 -4401
rect 19 -4435 31 -4401
rect -31 -4441 31 -4435
rect -125 -4503 125 -4497
rect -125 -4537 -113 -4503
rect 113 -4537 125 -4503
rect -125 -4543 125 -4537
<< properties >>
string FIXED_BBOX -178 -4520 178 4520
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 10.0 l 0.35 m 4 nf 1 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
