magic
tech sky130A
magscale 1 2
timestamp 1730482424
<< pwell >>
rect -1825 -2210 1825 2210
<< nmoslvt >>
rect -1629 -2000 -29 2000
rect 29 -2000 1629 2000
<< ndiff >>
rect -1687 1392 -1629 2000
rect -1687 -1392 -1675 1392
rect -1641 -1392 -1629 1392
rect -1687 -2000 -1629 -1392
rect -29 1392 29 2000
rect -29 -1392 -17 1392
rect 17 -1392 29 1392
rect -29 -2000 29 -1392
rect 1629 1392 1687 2000
rect 1629 -1392 1641 1392
rect 1675 -1392 1687 1392
rect 1629 -2000 1687 -1392
<< ndiffc >>
rect -1675 -1392 -1641 1392
rect -17 -1392 17 1392
rect 1641 -1392 1675 1392
<< psubdiff >>
rect -1789 2140 -1185 2174
rect 1185 2140 1789 2174
rect -1789 1455 -1755 2140
rect -1789 -2140 -1755 -1455
rect 1755 1455 1789 2140
rect 1755 -2140 1789 -1455
rect -1789 -2174 -1185 -2140
rect 1185 -2174 1789 -2140
<< psubdiffcont >>
rect -1185 2140 1185 2174
rect -1789 -1455 -1755 1455
rect 1755 -1455 1789 1455
rect -1185 -2174 1185 -2140
<< poly >>
rect -1394 2072 -264 2088
rect -1394 2055 -1378 2072
rect -1629 2038 -1378 2055
rect -280 2055 -264 2072
rect 264 2072 1394 2088
rect 264 2055 280 2072
rect -280 2038 -29 2055
rect -1629 2000 -29 2038
rect 29 2038 280 2055
rect 1378 2055 1394 2072
rect 1378 2038 1629 2055
rect 29 2000 1629 2038
rect -1629 -2038 -29 -2000
rect -1629 -2055 -1378 -2038
rect -1394 -2072 -1378 -2055
rect -280 -2055 -29 -2038
rect 29 -2038 1629 -2000
rect 29 -2055 280 -2038
rect -280 -2072 -264 -2055
rect -1394 -2088 -264 -2072
rect 264 -2072 280 -2055
rect 1378 -2055 1629 -2038
rect 1378 -2072 1394 -2055
rect 264 -2088 1394 -2072
<< polycont >>
rect -1378 2038 -280 2072
rect 280 2038 1378 2072
rect -1378 -2072 -280 -2038
rect 280 -2072 1378 -2038
<< locali >>
rect -1789 2140 -1229 2174
rect 1229 2140 1789 2174
rect -1789 1498 -1755 2140
rect 1755 1498 1789 2140
rect -1675 1392 -1641 1408
rect -1675 -1408 -1641 -1392
rect -17 1392 17 1408
rect -17 -1408 17 -1392
rect 1641 1392 1675 1408
rect 1641 -1408 1675 -1392
rect -1789 -2140 -1755 -1498
rect 1755 -2140 1789 -1498
rect -1789 -2174 -1229 -2140
rect 1229 -2174 1789 -2140
<< viali >>
rect -1229 2140 -1185 2174
rect -1185 2140 1185 2174
rect 1185 2140 1229 2174
rect -1613 2038 -1378 2072
rect -1378 2038 -280 2072
rect -280 2038 -45 2072
rect 45 2038 280 2072
rect 280 2038 1378 2072
rect 1378 2038 1613 2072
rect -1789 1455 -1755 1498
rect -1789 -1455 -1755 1455
rect 1755 1455 1789 1498
rect -1675 -1392 -1641 1392
rect -17 -1392 17 1392
rect 1641 -1392 1675 1392
rect -1789 -1498 -1755 -1455
rect 1755 -1455 1789 1455
rect 1755 -1498 1789 -1455
rect -1613 -2072 -1378 -2038
rect -1378 -2072 -280 -2038
rect -280 -2072 -45 -2038
rect 45 -2072 280 -2038
rect 280 -2072 1378 -2038
rect 1378 -2072 1613 -2038
rect -1229 -2174 -1185 -2140
rect -1185 -2174 1185 -2140
rect 1185 -2174 1229 -2140
<< metal1 >>
rect -1241 2174 1241 2180
rect -1241 2140 -1229 2174
rect 1229 2140 1241 2174
rect -1241 2134 1241 2140
rect -1625 2072 -33 2078
rect -1625 2038 -1613 2072
rect -45 2038 -33 2072
rect -1625 2032 -33 2038
rect 33 2072 1625 2078
rect 33 2038 45 2072
rect 1613 2038 1625 2072
rect 33 2032 1625 2038
rect -1795 1498 -1749 1510
rect -1795 -1498 -1789 1498
rect -1755 -1498 -1749 1498
rect 1749 1498 1795 1510
rect -1681 1392 -1635 1404
rect -1681 -1392 -1675 1392
rect -1641 -1392 -1635 1392
rect -1681 -1404 -1635 -1392
rect -23 1392 23 1404
rect -23 -1392 -17 1392
rect 17 -1392 23 1392
rect -23 -1404 23 -1392
rect 1635 1392 1681 1404
rect 1635 -1392 1641 1392
rect 1675 -1392 1681 1392
rect 1635 -1404 1681 -1392
rect -1795 -1510 -1749 -1498
rect 1749 -1498 1755 1498
rect 1789 -1498 1795 1498
rect 1749 -1510 1795 -1498
rect -1625 -2038 -33 -2032
rect -1625 -2072 -1613 -2038
rect -45 -2072 -33 -2038
rect -1625 -2078 -33 -2072
rect 33 -2038 1625 -2032
rect 33 -2072 45 -2038
rect 1613 -2072 1625 -2038
rect 33 -2078 1625 -2072
rect -1241 -2140 1241 -2134
rect -1241 -2174 -1229 -2140
rect 1229 -2174 1241 -2140
rect -1241 -2180 1241 -2174
<< properties >>
string FIXED_BBOX -1772 -2157 1772 2157
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 20.0 l 8.0 m 1 nf 2 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 70 viadrn 70 viagate 100 viagb 70 viagr 70 viagl 70 viagt 70
<< end >>
